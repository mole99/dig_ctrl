* NGSPICE file created from dig_ctrl_top.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlclkp_1 abstract view
.subckt sky130_fd_sc_hd__dlclkp_1 CLK GATE VGND VNB VPB VPWR GCLK
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlxtp_1 abstract view
.subckt sky130_fd_sc_hd__dlxtp_1 D GATE VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_4 abstract view
.subckt sky130_fd_sc_hd__o41a_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VPWR VGND VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_2 abstract view
.subckt sky130_fd_sc_hd__nor4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_4 abstract view
.subckt sky130_fd_sc_hd__or4b_4 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_2 abstract view
.subckt sky130_fd_sc_hd__o22a_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd1_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd1_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s4s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s4s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_4 abstract view
.subckt sky130_fd_sc_hd__nand4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_2 abstract view
.subckt sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_4 abstract view
.subckt sky130_fd_sc_hd__o211a_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_2 abstract view
.subckt sky130_fd_sc_hd__a2111oi_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_8 abstract view
.subckt sky130_fd_sc_hd__inv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_4 abstract view
.subckt sky130_fd_sc_hd__o22a_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlxtn_1 abstract view
.subckt sky130_fd_sc_hd__dlxtn_1 D GATE_N VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_2 abstract view
.subckt sky130_fd_sc_hd__nor3b_2 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_16 abstract view
.subckt sky130_fd_sc_hd__inv_16 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_4 abstract view
.subckt sky130_fd_sc_hd__o32a_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_12 abstract view
.subckt sky130_fd_sc_hd__inv_12 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_8 abstract view
.subckt sky130_fd_sc_hd__clkinv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_2 abstract view
.subckt sky130_fd_sc_hd__o41a_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_2 abstract view
.subckt sky130_fd_sc_hd__a22oi_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__bufinv_16 abstract view
.subckt sky130_fd_sc_hd__bufinv_16 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_1 abstract view
.subckt sky130_fd_sc_hd__a2111oi_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_6 abstract view
.subckt sky130_fd_sc_hd__inv_6 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_16 abstract view
.subckt sky130_fd_sc_hd__clkinv_16 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32ai_4 abstract view
.subckt sky130_fd_sc_hd__o32ai_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41ai_2 abstract view
.subckt sky130_fd_sc_hd__o41ai_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_2 abstract view
.subckt sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_4 abstract view
.subckt sky130_fd_sc_hd__o221ai_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_4 abstract view
.subckt sky130_fd_sc_hd__a221oi_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_4 abstract view
.subckt sky130_fd_sc_hd__and4bb_4 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_4 abstract view
.subckt sky130_fd_sc_hd__and4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_1 abstract view
.subckt sky130_fd_sc_hd__o221ai_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlxtn_2 abstract view
.subckt sky130_fd_sc_hd__dlxtn_2 D GATE_N VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41ai_4 abstract view
.subckt sky130_fd_sc_hd__o41ai_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_1 abstract view
.subckt sky130_fd_sc_hd__o2111ai_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_4 abstract view
.subckt sky130_fd_sc_hd__and3b_4 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_4 abstract view
.subckt sky130_fd_sc_hd__nor3b_4 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_4 abstract view
.subckt sky130_fd_sc_hd__a2111oi_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

.subckt dig_ctrl_top VDPWR VGND clk clk_o ena port_ms_i port_ms_o[0] port_ms_o[1]
+ port_ms_o[2] port_ms_o[3] port_ms_o[4] port_ms_o[5] port_ms_o[6] port_ms_o[7] rst_n
+ ui_in[0] ui_in[1] ui_in[2] ui_in[3] ui_in[4] ui_in[5] ui_in[6] ui_in[7] uio_in[0]
+ uio_in[1] uio_in[2] uio_in[3] uio_in[4] uio_in[5] uio_in[6] uio_in[7] uio_oe[0]
+ uio_oe[1] uio_oe[2] uio_oe[3] uio_oe[4] uio_oe[5] uio_oe[6] uio_oe[7] uio_out[0]
+ uio_out[1] uio_out[2] uio_out[3] uio_out[4] uio_out[5] uio_out[6] uio_out[7] uo_out[0]
+ uo_out[1] uo_out[2] uo_out[3] uo_out[4] uo_out[5] uo_out[6] uo_out[7]
X_2037_ _1010_ _0200_ VGND VGND VDPWR VDPWR _0741_ sky130_fd_sc_hd__and2_2
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[46\].clock_gate clknet_leaf_16_clk dig_ctrl_inst.latch_mem_inst.data_we\[46\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.gen_gclk\[46\]._gclk sky130_fd_sc_hd__dlclkp_1
X_2106_ dig_ctrl_inst.cpu_inst.data\[5\] dig_ctrl_inst.cpu_inst.data\[4\] dig_ctrl_inst.cpu_inst.data\[7\]
+ dig_ctrl_inst.cpu_inst.data\[6\] VGND VGND VDPWR VDPWR _0799_ sky130_fd_sc_hd__or4_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[41\].gen_latches\[3\].p_latch net221 dig_ctrl_inst.latch_mem_inst.gclk\[41\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[41\]\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_43_70 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_15_Left_93 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[30\].gen_latches\[1\].p_latch net234 dig_ctrl_inst.latch_mem_inst.gclk\[30\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[30\]\[1\] sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_68_570 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_470 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer7 _1079_ VGND VGND VDPWR VDPWR net289 sky130_fd_sc_hd__buf_2
XFILLER_0_64_14 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_6
X_1270_ _1018_ _1116_ _1115_ _1114_ _1117_ VGND VGND VDPWR VDPWR _1118_ sky130_fd_sc_hd__o41a_4
XFILLER_0_58_188 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[56\].gen_latches\[6\].p_latch net196 dig_ctrl_inst.latch_mem_inst.gclk\[56\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[56\]\[6\] sky130_fd_sc_hd__dlxtp_1
X_1606_ _0314_ _0315_ _0316_ _0317_ VGND VGND VDPWR VDPWR _0318_ sky130_fd_sc_hd__or4_1
XFILLER_0_14_203 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_1468_ _0194_ _0196_ VGND VGND VDPWR VDPWR _0009_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_57_507 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout127 _1128_ VGND VGND VDPWR VDPWR net127 sky130_fd_sc_hd__clkbuf_2
Xfanout138 _0227_ VGND VGND VDPWR VDPWR net138 sky130_fd_sc_hd__buf_2
Xfanout105 _1134_ VGND VGND VDPWR VDPWR net105 sky130_fd_sc_hd__buf_4
X_1399_ net148 _0154_ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.data_we\[57\]
+ sky130_fd_sc_hd__and2_1
Xfanout149 net151 VGND VGND VDPWR VDPWR net149 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout116 net117 VGND VGND VDPWR VDPWR net116 sky130_fd_sc_hd__buf_4
X_1537_ net171 net169 VGND VGND VDPWR VDPWR _0250_ sky130_fd_sc_hd__nor2_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[45\].gen_latches\[4\].p_latch net210 dig_ctrl_inst.latch_mem_inst.gclk\[45\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[45\]\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_64_125 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_309 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_40_407 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[34\].gen_latches\[2\].p_latch net227 dig_ctrl_inst.latch_mem_inst.gclk\[34\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[34\]\[2\] sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_0_Left_78 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_5_195 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_29 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[23\].gen_latches\[0\].p_latch net247 dig_ctrl_inst.latch_mem_inst.gclk\[23\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[23\]\[0\] sky130_fd_sc_hd__dlxtp_1
X_2440_ clknet_leaf_6_clk _0048_ net145 VGND VGND VDPWR VDPWR dig_ctrl_inst.cpu_inst.r0\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_55_169 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_320 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_69 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
X_1253_ net257 dig_ctrl_inst.cpu_inst.r1\[5\] VGND VGND VDPWR VDPWR _1101_ sky130_fd_sc_hd__and2b_1
X_2371_ net248 _0990_ _0995_ _0997_ VGND VGND VDPWR VDPWR _0111_ sky130_fd_sc_hd__a22o_1
X_1322_ net129 net66 VGND VGND VDPWR VDPWR _0119_ sky130_fd_sc_hd__and2_1
X_1184_ net260 net256 dig_ctrl_inst.cpu_inst.r3\[3\] VGND VGND VDPWR VDPWR _1032_
+ sky130_fd_sc_hd__and3_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[11\].gen_latches\[7\].p_latch net188 dig_ctrl_inst.latch_mem_inst.gclk\[11\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[11\]\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_46_136 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_233 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[5\].gen_latches\[0\].p_latch net243 dig_ctrl_inst.latch_mem_inst.gclk\[5\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[5\]\[0\] sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_27_Left_105 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[49\].gen_latches\[5\].p_latch net199 dig_ctrl_inst.latch_mem_inst.gclk\[49\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[49\]\[5\] sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_2_176 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_36_Left_114 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[38\].gen_latches\[3\].p_latch net216 dig_ctrl_inst.latch_mem_inst.gclk\[38\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[38\]\[3\] sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[27\].gen_latches\[1\].p_latch net237 dig_ctrl_inst.latch_mem_inst.gclk\[27\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[27\]\[1\] sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_45_Left_123 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_29 VDPWR VGND VDPWR VGND sky130_ef_sc_hd__decap_12
X_1940_ dig_ctrl_inst.latch_mem_inst.RAM\[30\]\[6\] net74 net70 VGND VGND VDPWR VDPWR
+ _0646_ sky130_fd_sc_hd__and3_2
X_1871_ _0577_ _0568_ _0570_ _0287_ VGND VGND VDPWR VDPWR _0578_ sky130_fd_sc_hd__nor4_2
XPHY_EDGE_ROW_54_Left_132 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_139 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_309 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_85 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
X_2423_ clknet_leaf_13_clk _0031_ net139 VGND VGND VDPWR VDPWR dig_ctrl_inst.cpu_inst.instr\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_2354_ dig_ctrl_inst.cpu_inst.port_o\[0\] net17 _0988_ VGND VGND VDPWR VDPWR _0103_
+ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_63_Left_141 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
X_1236_ _1018_ _1082_ _1081_ _1080_ _1083_ VGND VGND VDPWR VDPWR _1084_ sky130_fd_sc_hd__o41a_4
X_2285_ _0752_ _0830_ _0833_ VGND VGND VDPWR VDPWR _0969_ sky130_fd_sc_hd__a21o_1
X_1305_ net150 _1143_ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.data_we\[9\]
+ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_72_Left_150 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
X_1167_ dig_ctrl_inst.cpu_inst.instr\[7\] dig_ctrl_inst.cpu_inst.instr\[6\] net252
+ net253 VGND VGND VDPWR VDPWR _1015_ sky130_fd_sc_hd__or4b_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[9\].gen_latches\[1\].p_latch net232 dig_ctrl_inst.latch_mem_inst.gclk\[9\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[9\]\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_19_169 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_73_605 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_392 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_292 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_334 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
X_2070_ _0761_ _0762_ _1068_ VGND VGND VDPWR VDPWR _0763_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_3_Left_81 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_328 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_223 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_1854_ dig_ctrl_inst.latch_mem_inst.RAM\[13\]\[4\] _0114_ _0129_ dig_ctrl_inst.latch_mem_inst.RAM\[26\]\[4\]
+ VGND VGND VDPWR VDPWR _0562_ sky130_fd_sc_hd__a22o_1
X_1923_ dig_ctrl_inst.latch_mem_inst.RAM\[2\]\[6\] net121 net112 VGND VGND VDPWR VDPWR
+ _0629_ sky130_fd_sc_hd__and3_2
X_1785_ dig_ctrl_inst.latch_mem_inst.RAM\[33\]\[3\] _0135_ _0491_ _0492_ _0493_ VGND
+ VGND VDPWR VDPWR _0494_ sky130_fd_sc_hd__a2111o_1
X_2406_ clknet_leaf_5_clk _0014_ net146 VGND VGND VDPWR VDPWR dig_ctrl_inst.cpu_inst.port_o\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_183 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_194 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
X_2337_ dig_ctrl_inst.cpu_inst.port_o\[1\] net357 _0986_ VGND VGND VDPWR VDPWR _0088_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_3 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_27_329 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1219_ dig_ctrl_inst.cpu_inst.r0\[0\] _1019_ _1065_ _1066_ VGND VGND VDPWR VDPWR
+ _1067_ sky130_fd_sc_hd__o22a_2
X_2268_ _0836_ _0908_ _0953_ VGND VGND VDPWR VDPWR _0954_ sky130_fd_sc_hd__o21a_1
X_2199_ _0836_ _0837_ _0887_ _0770_ _0886_ VGND VGND VDPWR VDPWR _0888_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_35_373 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_150 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[53\].clock_gate clknet_leaf_17_clk dig_ctrl_inst.latch_mem_inst.data_we\[53\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.gen_gclk\[53\]._gclk sky130_fd_sc_hd__dlclkp_1
XFILLER_0_22_109 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_6
Xhold63 dig_ctrl_inst.spi_receiver_inst.spi_mosi_sync VGND VGND VDPWR VDPWR net345
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold52 dig_ctrl_inst.synchronizer_port_i_inst\[2\].pipe\[0\] VGND VGND VDPWR VDPWR
+ net334 sky130_fd_sc_hd__dlygate4sd3_1
Xhold74 dig_ctrl_inst.spi_data_i\[5\] VGND VGND VDPWR VDPWR net356 sky130_fd_sc_hd__dlygate4sd3_1
Xhold41 dig_ctrl_inst.latch_mem_inst.wdata\[4\] VGND VGND VDPWR VDPWR net323 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_29 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
Xhold96 dig_ctrl_inst.cpu_inst.r2\[4\] VGND VGND VDPWR VDPWR net378 sky130_fd_sc_hd__dlygate4sd3_1
Xhold85 dig_ctrl_inst.cpu_inst.r1\[1\] VGND VGND VDPWR VDPWR net367 sky130_fd_sc_hd__dlygate4sd3_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[60\].gen_latches\[1\].p_latch net234 dig_ctrl_inst.latch_mem_inst.gclk\[60\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[60\]\[1\] sky130_fd_sc_hd__dlxtp_1
X_1570_ net123 net119 net82 net68 net130 VGND VGND VDPWR VDPWR _0282_ sky130_fd_sc_hd__a32o_1
XANTENNA_5 _0560_ VGND VGND VDPWR VDPWR sky130_fd_sc_hd__diode_2
XFILLER_0_21_164 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
Xrebuffer17 net300 VGND VGND VDPWR VDPWR net299 sky130_fd_sc_hd__dlygate4sd1_1
X_2122_ net157 net138 net137 VGND VGND VDPWR VDPWR _0814_ sky130_fd_sc_hd__and3_2
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[52\].clock_buffer dig_ctrl_inst.latch_mem_inst.gen_gclk\[52\]._gclk
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.gclk\[52\] sky130_fd_sc_hd__clkbuf_4
X_2053_ net254 _1015_ _0744_ _0745_ VGND VGND VDPWR VDPWR _0746_ sky130_fd_sc_hd__o211a_1
XFILLER_0_44_201 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_32_354 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_73 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_2528__275 VGND VGND VDPWR VDPWR _2528__275/HI net275 sky130_fd_sc_hd__conb_1
X_1837_ dig_ctrl_inst.latch_mem_inst.RAM\[43\]\[4\] net108 net92 net58 VGND VGND VDPWR
+ VDPWR _0545_ sky130_fd_sc_hd__and4_1
X_1906_ dig_ctrl_inst.latch_mem_inst.RAM\[44\]\[5\] net76 net52 VGND VGND VDPWR VDPWR
+ _0613_ sky130_fd_sc_hd__and3_2
X_1768_ dig_ctrl_inst.latch_mem_inst.RAM\[55\]\[3\] _0153_ _0474_ _0475_ _0476_ VGND
+ VGND VDPWR VDPWR _0477_ sky130_fd_sc_hd__a2111o_1
X_1699_ dig_ctrl_inst.latch_mem_inst.RAM\[10\]\[2\] net126 net85 VGND VGND VDPWR VDPWR
+ _0409_ sky130_fd_sc_hd__and3_2
XFILLER_0_12_197 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_337 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
Xoutput31 net31 VGND VGND VDPWR VDPWR uo_out[3] sky130_fd_sc_hd__buf_2
Xoutput20 net20 VGND VGND VDPWR VDPWR port_ms_o[3] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_54_490 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[53\].gen_latches\[0\].p_latch net242 dig_ctrl_inst.latch_mem_inst.gclk\[53\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[53\]\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_26_201 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_1622_ dig_ctrl_inst.latch_mem_inst.RAM\[9\]\[0\] _1143_ _0295_ _0299_ _0304_ VGND
+ VGND VDPWR VDPWR _0334_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_1_301 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_1484_ dig_ctrl_inst.cpu_inst.skip _0173_ _0202_ VGND VGND VDPWR VDPWR _0203_ sky130_fd_sc_hd__a21o_1
X_1553_ net166 _0252_ net167 VGND VGND VDPWR VDPWR _0266_ sky130_fd_sc_hd__nand3b_1
X_2105_ _0782_ _0789_ _0796_ _0797_ VGND VGND VDPWR VDPWR _0798_ sky130_fd_sc_hd__and4_1
X_2036_ dig_ctrl_inst.cpu_inst.instr\[7\] _0740_ _0276_ VGND VGND VDPWR VDPWR _0033_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_72_340 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[41\].gen_latches\[7\].p_latch net184 dig_ctrl_inst.latch_mem_inst.gclk\[41\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[41\]\[7\] sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_68_571 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[30\].gen_latches\[5\].p_latch net205 dig_ctrl_inst.latch_mem_inst.gclk\[30\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[30\]\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_55_318 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
Xrebuffer8 net291 VGND VGND VDPWR VDPWR net290 sky130_fd_sc_hd__dlymetal6s4s_1
XTAP_TAPCELL_ROW_51_471 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_37 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[57\].gen_latches\[1\].p_latch net232 dig_ctrl_inst.latch_mem_inst.gclk\[57\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[57\]\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_13_30 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_1536_ net170 net169 VGND VGND VDPWR VDPWR _0249_ sky130_fd_sc_hd__nand2_1
X_1605_ dig_ctrl_inst.latch_mem_inst.RAM\[16\]\[0\] _0119_ _0137_ dig_ctrl_inst.latch_mem_inst.RAM\[35\]\[0\]
+ VGND VGND VDPWR VDPWR _0317_ sky130_fd_sc_hd__a22o_1
Xfanout106 net107 VGND VGND VDPWR VDPWR net106 sky130_fd_sc_hd__buf_4
X_1467_ _1096_ _0195_ _0184_ VGND VGND VDPWR VDPWR _0196_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_57_508 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_60 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_8
Xfanout139 net140 VGND VGND VDPWR VDPWR net139 sky130_fd_sc_hd__clkbuf_4
Xfanout117 _1129_ VGND VGND VDPWR VDPWR net117 sky130_fd_sc_hd__buf_4
X_1398_ net114 net90 net42 VGND VGND VDPWR VDPWR _0154_ sky130_fd_sc_hd__and3_4
Xfanout128 net130 VGND VGND VDPWR VDPWR net128 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_65_552 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2019_ dig_ctrl_inst.latch_mem_inst.RAM\[3\]\[7\] _1135_ _0120_ dig_ctrl_inst.latch_mem_inst.RAM\[17\]\[7\]
+ _0723_ VGND VGND VDPWR VDPWR _0724_ sky130_fd_sc_hd__a221o_1
XFILLER_0_54_81 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[1\].gen_latches\[3\].p_latch net220 dig_ctrl_inst.latch_mem_inst.gclk\[1\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[1\]\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_9_231 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[34\].gen_latches\[6\].p_latch net191 dig_ctrl_inst.latch_mem_inst.gclk\[34\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[34\]\[6\] sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_5_196 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_588 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_17 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[23\].gen_latches\[4\].p_latch net211 dig_ctrl_inst.latch_mem_inst.gclk\[23\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[23\]\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_59_48 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_8
Xdig_ctrl_inst.latch_mem_inst.gen_words\[12\].gen_latches\[2\].p_latch net231 dig_ctrl_inst.latch_mem_inst.gclk\[12\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[12\]\[2\] sky130_fd_sc_hd__dlxtp_1
X_1321_ _1112_ _1127_ VGND VGND VDPWR VDPWR _0118_ sky130_fd_sc_hd__and2b_1
X_1252_ net261 net257 dig_ctrl_inst.cpu_inst.r3\[5\] VGND VGND VDPWR VDPWR _1100_
+ sky130_fd_sc_hd__and3_2
X_2370_ _0990_ _0996_ VGND VGND VDPWR VDPWR _0997_ sky130_fd_sc_hd__nor2_1
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[45\].clock_buffer dig_ctrl_inst.latch_mem_inst.gen_gclk\[45\]._gclk
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.gclk\[45\] sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_19_276 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_73 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
X_1183_ net258 net254 VGND VGND VDPWR VDPWR _1031_ sky130_fd_sc_hd__nand2_1
XFILLER_0_40_83 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_2499_ clknet_leaf_5_clk _0096_ net177 VGND VGND VDPWR VDPWR net29 sky130_fd_sc_hd__dfrtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[58\].clock_gate clknet_leaf_1_clk dig_ctrl_inst.latch_mem_inst.data_we\[58\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.gen_gclk\[58\]._gclk sky130_fd_sc_hd__dlclkp_1
XFILLER_0_64_3 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
X_1519_ _0998_ dig_ctrl_inst.cpu_inst.r2\[7\] dig_ctrl_inst.cpu_inst.r1\[7\] _1022_
+ net299 VGND VGND VDPWR VDPWR _0232_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_12_Right_12 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[5\].gen_latches\[4\].p_latch net213 dig_ctrl_inst.latch_mem_inst.gclk\[5\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[5\]\[4\] sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_2_177 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_21_Right_21 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_148 VDPWR VGND VDPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_181 VDPWR VGND VDPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_30_Right_30 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[38\].gen_latches\[7\].p_latch net184 dig_ctrl_inst.latch_mem_inst.gclk\[38\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[38\]\[7\] sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[60\].clock_gate clknet_leaf_0_clk dig_ctrl_inst.latch_mem_inst.data_we\[60\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.gen_gclk\[60\]._gclk sky130_fd_sc_hd__dlclkp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[27\].gen_latches\[5\].p_latch net204 dig_ctrl_inst.latch_mem_inst.gclk\[27\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[27\]\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_28_115 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_1870_ _0574_ _0575_ _0576_ VGND VGND VDPWR VDPWR _0577_ sky130_fd_sc_hd__or3_1
XFILLER_0_36_181 VDPWR VGND VDPWR VGND sky130_ef_sc_hd__decap_12
X_2353_ dig_ctrl_inst.cpu_inst.data\[0\] dig_ctrl_inst.cpu_inst.port_stb_o _0800_
+ _0801_ VGND VGND VDPWR VDPWR _0988_ sky130_fd_sc_hd__nand4_4
X_2422_ clknet_leaf_13_clk _0030_ net139 VGND VGND VDPWR VDPWR dig_ctrl_inst.cpu_inst.instr\[4\]
+ sky130_fd_sc_hd__dfrtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[16\].gen_latches\[3\].p_latch net217 dig_ctrl_inst.latch_mem_inst.gclk\[16\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[16\]\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_35_61 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_1235_ net259 net255 dig_ctrl_inst.cpu_inst.r0\[1\] VGND VGND VDPWR VDPWR _1083_
+ sky130_fd_sc_hd__or3_1
X_2284_ net374 _0968_ _0967_ VGND VGND VDPWR VDPWR _0053_ sky130_fd_sc_hd__mux2_1
X_1304_ net120 net116 net90 VGND VGND VDPWR VDPWR _1143_ sky130_fd_sc_hd__and3_4
X_1166_ net252 net253 VGND VGND VDPWR VDPWR _1014_ sky130_fd_sc_hd__nand2b_1
X_1999_ dig_ctrl_inst.latch_mem_inst.RAM\[48\]\[7\] net129 net43 VGND VGND VDPWR VDPWR
+ _0704_ sky130_fd_sc_hd__and3_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[9\].gen_latches\[5\].p_latch net200 dig_ctrl_inst.latch_mem_inst.gclk\[9\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[9\]\[5\] sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_38_393 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[2\].clock_buffer dig_ctrl_inst.latch_mem_inst.gen_gclk\[2\]._gclk
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.gclk\[2\] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_33_195 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_21_293 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_27 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_1922_ dig_ctrl_inst.latch_mem_inst.RAM\[48\]\[6\] net129 net43 VGND VGND VDPWR VDPWR
+ _0628_ sky130_fd_sc_hd__and3_2
X_1853_ dig_ctrl_inst.latch_mem_inst.RAM\[21\]\[4\] _0124_ _0135_ dig_ctrl_inst.latch_mem_inst.RAM\[33\]\[4\]
+ VGND VGND VDPWR VDPWR _0561_ sky130_fd_sc_hd__a22o_1
X_1784_ dig_ctrl_inst.latch_mem_inst.RAM\[23\]\[3\] net103 net99 net62 VGND VGND VDPWR
+ VDPWR _0493_ sky130_fd_sc_hd__and4_1
XFILLER_0_12_324 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_63 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_2336_ dig_ctrl_inst.cpu_inst.port_o\[0\] net380 _0986_ VGND VGND VDPWR VDPWR _0087_
+ sky130_fd_sc_hd__mux2_1
X_2405_ clknet_leaf_6_clk _0013_ net146 VGND VGND VDPWR VDPWR dig_ctrl_inst.cpu_inst.port_o\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_1149_ net265 VGND VGND VDPWR VDPWR _0998_ sky130_fd_sc_hd__inv_2
X_1218_ net258 dig_ctrl_inst.cpu_inst.r2\[0\] VGND VGND VDPWR VDPWR _1066_ sky130_fd_sc_hd__and2b_1
X_2198_ _0761_ _0776_ _1068_ VGND VGND VDPWR VDPWR _0887_ sky130_fd_sc_hd__mux2_1
X_2267_ _0768_ _0817_ _0952_ _0770_ _0886_ VGND VGND VDPWR VDPWR _0953_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_35_374 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_165 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
Xhold53 dig_ctrl_inst.synchronizer_mode_i_inst.pipe\[0\] VGND VGND VDPWR VDPWR net335
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold75 dig_ctrl_inst.spi_data_i\[1\] VGND VGND VDPWR VDPWR net357 sky130_fd_sc_hd__dlygate4sd3_1
Xhold42 dig_ctrl_inst.latch_mem_inst.wdata\[2\] VGND VGND VDPWR VDPWR net324 sky130_fd_sc_hd__dlygate4sd3_1
Xhold64 dig_ctrl_inst.cpu_inst.prev_state\[0\] VGND VGND VDPWR VDPWR net346 sky130_fd_sc_hd__dlygate4sd3_1
Xhold86 dig_ctrl_inst.cpu_inst.r3\[5\] VGND VGND VDPWR VDPWR net368 sky130_fd_sc_hd__dlygate4sd3_1
Xhold97 dig_ctrl_inst.cpu_inst.r2\[0\] VGND VGND VDPWR VDPWR net379 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_232 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[60\].gen_latches\[5\].p_latch net203 dig_ctrl_inst.latch_mem_inst.gclk\[60\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[60\]\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_53_279 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XANTENNA_6 _0592_ VGND VGND VDPWR VDPWR sky130_fd_sc_hd__diode_2
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[38\].clock_buffer dig_ctrl_inst.latch_mem_inst.gen_gclk\[38\]._gclk
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.gclk\[38\] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_21_154 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
X_2121_ _0772_ _0810_ _0812_ VGND VGND VDPWR VDPWR _0813_ sky130_fd_sc_hd__and3_2
XFILLER_0_16_41 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
X_2052_ dig_ctrl_inst.cpu_inst.instr\[7\] dig_ctrl_inst.cpu_inst.instr\[6\] VGND VGND
+ VDPWR VDPWR _0745_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_76_338 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_32_355 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_95 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
X_1905_ dig_ctrl_inst.latch_mem_inst.RAM\[22\]\[5\] net93 net61 VGND VGND VDPWR VDPWR
+ _0612_ sky130_fd_sc_hd__and3_2
X_1836_ dig_ctrl_inst.latch_mem_inst.RAM\[14\]\[4\] net123 net72 VGND VGND VDPWR VDPWR
+ _0544_ sky130_fd_sc_hd__and3_2
X_1698_ dig_ctrl_inst.latch_mem_inst.RAM\[8\]\[2\] net122 net87 VGND VGND VDPWR VDPWR
+ _0408_ sky130_fd_sc_hd__and3_2
XPHY_EDGE_ROW_6_Right_6 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
X_1767_ dig_ctrl_inst.latch_mem_inst.RAM\[35\]\[3\] net131 net102 net51 VGND VGND
+ VDPWR VDPWR _0476_ sky130_fd_sc_hd__and4_1
X_2319_ dig_ctrl_inst.spi_data_i\[3\] dig_ctrl_inst.spi_data_i\[2\] dig_ctrl_inst.spi_receiver_inst.spi_cnt\[0\]
+ VGND VGND VDPWR VDPWR _0980_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_23_300 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput32 net32 VGND VGND VDPWR VDPWR uo_out[4] sky130_fd_sc_hd__buf_2
Xoutput21 net21 VGND VGND VDPWR VDPWR port_ms_o[4] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_59_Right_59 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_54_491 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_335 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_1552_ _0257_ _0264_ _0263_ VGND VGND VDPWR VDPWR _0265_ sky130_fd_sc_hd__a21oi_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[53\].gen_latches\[4\].p_latch net208 dig_ctrl_inst.latch_mem_inst.gclk\[53\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[53\]\[4\] sky130_fd_sc_hd__dlxtp_1
X_1621_ dig_ctrl_inst.latch_mem_inst.RAM\[41\]\[0\] _0141_ _0292_ _0298_ _0303_ VGND
+ VGND VDPWR VDPWR _0333_ sky130_fd_sc_hd__a2111o_1
XPHY_EDGE_ROW_68_Right_68 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
X_1483_ net248 dig_ctrl_inst.cpu_inst.cpu_state\[1\] _0999_ VGND VGND VDPWR VDPWR
+ _0202_ sky130_fd_sc_hd__o21ai_1
X_2104_ _0259_ _0785_ _0793_ _0258_ _0795_ VGND VGND VDPWR VDPWR _0797_ sky130_fd_sc_hd__o221a_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[42\].gen_latches\[2\].p_latch net230 dig_ctrl_inst.latch_mem_inst.gclk\[42\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[42\]\[2\] sky130_fd_sc_hd__dlxtp_1
X_2035_ _0728_ _0739_ _0729_ _0686_ VGND VGND VDPWR VDPWR _0740_ sky130_fd_sc_hd__o31a_1
XPHY_EDGE_ROW_77_Right_77 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_213 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_8
Xdig_ctrl_inst.latch_mem_inst.gen_words\[31\].gen_latches\[0\].p_latch net246 dig_ctrl_inst.latch_mem_inst.gclk\[31\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[31\]\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_25_290 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_162 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_50 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_6
X_1819_ dig_ctrl_inst.latch_mem_inst.RAM\[53\]\[4\] _0151_ _0524_ _0525_ _0526_ VGND
+ VGND VDPWR VDPWR _0527_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_68_572 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_113 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_51_472 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer9 net302 VGND VGND VDPWR VDPWR net291 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_16_290 VDPWR VGND VDPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_27 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_17 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_19 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[57\].gen_latches\[5\].p_latch net202 dig_ctrl_inst.latch_mem_inst.gclk\[57\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[57\]\[5\] sky130_fd_sc_hd__dlxtp_1
Xfanout107 net108 VGND VGND VDPWR VDPWR net107 sky130_fd_sc_hd__buf_4
Xfanout118 net119 VGND VGND VDPWR VDPWR net118 sky130_fd_sc_hd__clkbuf_2
X_1604_ dig_ctrl_inst.latch_mem_inst.RAM\[36\]\[0\] net98 net59 _0114_ dig_ctrl_inst.latch_mem_inst.RAM\[13\]\[0\]
+ VGND VGND VDPWR VDPWR _0316_ sky130_fd_sc_hd__a32o_1
Xfanout129 net130 VGND VGND VDPWR VDPWR net129 sky130_fd_sc_hd__clkbuf_2
X_1535_ _0246_ _0247_ VGND VGND VDPWR VDPWR _0248_ sky130_fd_sc_hd__nand2_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[46\].gen_latches\[3\].p_latch net217 dig_ctrl_inst.latch_mem_inst.gclk\[46\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[46\]\[3\] sky130_fd_sc_hd__dlxtp_1
X_1397_ net153 net88 net48 VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.data_we\[56\]
+ sky130_fd_sc_hd__and3_2
X_1466_ dig_ctrl_inst.spi_addr\[3\] dig_ctrl_inst.spi_addr\[4\] _0191_ VGND VGND VDPWR
+ VDPWR _0195_ sky130_fd_sc_hd__nand3_1
XTAP_TAPCELL_ROW_57_509 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_553 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2018_ dig_ctrl_inst.latch_mem_inst.RAM\[32\]\[7\] _0134_ _0279_ dig_ctrl_inst.latch_mem_inst.RAM\[6\]\[7\]
+ VGND VGND VDPWR VDPWR _0723_ sky130_fd_sc_hd__a22o_1
XFILLER_0_54_93 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[35\].gen_latches\[1\].p_latch net235 dig_ctrl_inst.latch_mem_inst.gclk\[35\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[35\]\[1\] sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[1\].gen_latches\[7\].p_latch net185 dig_ctrl_inst.latch_mem_inst.gclk\[1\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[1\]\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_9_287 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_260 VDPWR VGND VDPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_197 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_589 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1320_ net155 _0117_ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.data_we\[15\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_59_16 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_1251_ net260 net257 dig_ctrl_inst.cpu_inst.r2\[5\] VGND VGND VDPWR VDPWR _1099_
+ sky130_fd_sc_hd__and3b_1
X_1182_ _1025_ _1010_ VGND VGND VDPWR VDPWR _1030_ sky130_fd_sc_hd__and2_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[12\].gen_latches\[6\].p_latch net191 dig_ctrl_inst.latch_mem_inst.gclk\[12\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[12\]\[6\] sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_62_534 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_277 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_85 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
XFILLER_0_40_73 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_341 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_2498_ clknet_leaf_5_clk _0095_ net177 VGND VGND VDPWR VDPWR net28 sky130_fd_sc_hd__dfrtp_1
X_1449_ _0182_ _0183_ VGND VGND VDPWR VDPWR _0003_ sky130_fd_sc_hd__nor2_1
XFILLER_0_57_3 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
X_1518_ net265 net262 dig_ctrl_inst.cpu_inst.r3\[7\] VGND VGND VDPWR VDPWR _0231_
+ sky130_fd_sc_hd__and3_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[39\].gen_latches\[2\].p_latch net231 dig_ctrl_inst.latch_mem_inst.gclk\[39\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[39\]\[2\] sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_2_178 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_193 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_290 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[28\].gen_latches\[0\].p_latch net240 dig_ctrl_inst.latch_mem_inst.gclk\[28\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[28\]\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_45_18 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_16_258 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_193 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
X_2352_ dig_ctrl_inst.cpu_inst.port_o\[7\] net35 _0987_ VGND VGND VDPWR VDPWR _0102_
+ sky130_fd_sc_hd__mux2_1
X_1303_ net155 net126 net89 VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.data_we\[8\]
+ sky130_fd_sc_hd__and3_2
X_2421_ clknet_leaf_9_clk _0029_ net141 VGND VGND VDPWR VDPWR dig_ctrl_inst.cpu_inst.arg1\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_2283_ net164 _0751_ _0798_ VGND VGND VDPWR VDPWR _0968_ sky130_fd_sc_hd__o21ai_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[16\].gen_latches\[7\].p_latch net184 dig_ctrl_inst.latch_mem_inst.gclk\[16\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[16\]\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_35_40 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
X_1234_ net255 dig_ctrl_inst.cpu_inst.r1\[1\] VGND VGND VDPWR VDPWR _1082_ sky130_fd_sc_hd__and2b_1
X_1165_ dig_ctrl_inst.cpu_inst.instr\[6\] dig_ctrl_inst.cpu_inst.instr\[7\] VGND VGND
+ VDPWR VDPWR _1013_ sky130_fd_sc_hd__nor2_1
XFILLER_0_27_160 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_8
X_1998_ dig_ctrl_inst.latch_mem_inst.RAM\[26\]\[7\] net83 net70 VGND VGND VDPWR VDPWR
+ _0703_ sky130_fd_sc_hd__and3_2
XFILLER_0_42_141 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_7_204 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_394 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire113 _1132_ VGND VGND VDPWR VDPWR net113 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_25_119 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_6
X_1852_ dig_ctrl_inst.latch_mem_inst.RAM\[15\]\[4\] _0117_ _0159_ dig_ctrl_inst.latch_mem_inst.RAM\[62\]\[4\]
+ VGND VGND VDPWR VDPWR _0560_ sky130_fd_sc_hd__a22o_1
X_1921_ dig_ctrl_inst.latch_mem_inst.RAM\[19\]\[6\] net133 net104 net66 VGND VGND
+ VDPWR VDPWR _0627_ sky130_fd_sc_hd__and4_1
XFILLER_0_16_108 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
X_1783_ dig_ctrl_inst.latch_mem_inst.RAM\[2\]\[3\] net122 net110 VGND VGND VDPWR VDPWR
+ _0492_ sky130_fd_sc_hd__and3_2
X_2335_ dig_ctrl_inst.cpu_inst.port_stb_o _0804_ VGND VGND VDPWR VDPWR _0986_ sky130_fd_sc_hd__nand2_4
X_2404_ clknet_leaf_6_clk _0012_ net146 VGND VGND VDPWR VDPWR dig_ctrl_inst.cpu_inst.port_o\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_2266_ _0814_ _0817_ VGND VGND VDPWR VDPWR _0952_ sky130_fd_sc_hd__and2b_1
XFILLER_0_46_83 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_1217_ dig_ctrl_inst.cpu_inst.r1\[0\] _1000_ _1018_ _1064_ VGND VGND VDPWR VDPWR
+ _1065_ sky130_fd_sc_hd__a211o_1
X_2197_ net168 _0769_ VGND VGND VDPWR VDPWR _0886_ sky130_fd_sc_hd__nand2_1
XFILLER_0_47_288 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_35_375 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_341 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_163 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[61\].gen_latches\[0\].p_latch net242 dig_ctrl_inst.latch_mem_inst.gclk\[61\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[61\]\[0\] sky130_fd_sc_hd__dlxtp_1
Xhold54 dig_ctrl_inst.spi_receiver_inst.synchronizer_spi_mosi.pipe\[0\] VGND VGND
+ VDPWR VDPWR net336 sky130_fd_sc_hd__dlygate4sd3_1
Xhold98 dig_ctrl_inst.spi_data_i\[0\] VGND VGND VDPWR VDPWR net380 sky130_fd_sc_hd__dlygate4sd3_1
Xhold87 dig_ctrl_inst.cpu_inst.r1\[2\] VGND VGND VDPWR VDPWR net369 sky130_fd_sc_hd__dlygate4sd3_1
Xhold43 dig_ctrl_inst.latch_mem_inst.wdata\[0\] VGND VGND VDPWR VDPWR net325 sky130_fd_sc_hd__dlygate4sd3_1
Xhold65 _0042_ VGND VGND VDPWR VDPWR net347 sky130_fd_sc_hd__dlygate4sd3_1
Xhold76 dig_ctrl_inst.cpu_inst.r3\[1\] VGND VGND VDPWR VDPWR net358 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_26_320 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_247 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XANTENNA_7 _0666_ VGND VGND VDPWR VDPWR sky130_fd_sc_hd__diode_2
X_2120_ _0765_ _0808_ _0811_ _0768_ VGND VGND VDPWR VDPWR _0812_ sky130_fd_sc_hd__o22a_1
Xrebuffer19 _1094_ VGND VGND VDPWR VDPWR net301 sky130_fd_sc_hd__dlygate4sd1_1
XTAP_TAPCELL_ROW_49_456 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2051_ dig_ctrl_inst.cpu_inst.instr\[6\] dig_ctrl_inst.cpu_inst.instr\[7\] VGND VGND
+ VDPWR VDPWR _0744_ sky130_fd_sc_hd__nand2b_2
X_1835_ dig_ctrl_inst.latch_mem_inst.RAM\[38\]\[4\] net95 net58 VGND VGND VDPWR VDPWR
+ _0543_ sky130_fd_sc_hd__and3_2
XTAP_TAPCELL_ROW_32_356 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1904_ dig_ctrl_inst.latch_mem_inst.RAM\[15\]\[5\] _0117_ _0608_ _0609_ _0610_ VGND
+ VGND VDPWR VDPWR _0611_ sky130_fd_sc_hd__a2111o_1
X_1697_ dig_ctrl_inst.latch_mem_inst.RAM\[20\]\[2\] net97 net71 VGND VGND VDPWR VDPWR
+ _0407_ sky130_fd_sc_hd__and3_2
X_1766_ dig_ctrl_inst.latch_mem_inst.RAM\[38\]\[3\] net93 net53 VGND VGND VDPWR VDPWR
+ _0475_ sky130_fd_sc_hd__and3_2
X_2318_ dig_ctrl_inst.spi_data_i\[7\] dig_ctrl_inst.spi_data_i\[6\] dig_ctrl_inst.spi_data_i\[5\]
+ dig_ctrl_inst.spi_data_i\[4\] dig_ctrl_inst.spi_receiver_inst.spi_cnt\[0\] dig_ctrl_inst.spi_receiver_inst.spi_cnt\[1\]
+ VGND VGND VDPWR VDPWR _0979_ sky130_fd_sc_hd__mux4_1
X_2249_ _0747_ _0749_ _0935_ VGND VGND VDPWR VDPWR _0936_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_23_301 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput33 net33 VGND VGND VDPWR VDPWR uo_out[5] sky130_fd_sc_hd__buf_2
Xoutput22 net22 VGND VGND VDPWR VDPWR port_ms_o[5] sky130_fd_sc_hd__buf_2
XFILLER_0_9_3 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_206 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
X_1482_ _0200_ _1027_ VGND VGND VDPWR VDPWR _0201_ sky130_fd_sc_hd__nand2b_1
X_1551_ _1068_ net164 VGND VGND VDPWR VDPWR _0264_ sky130_fd_sc_hd__nand2_1
X_1620_ dig_ctrl_inst.latch_mem_inst.RAM\[33\]\[0\] _0135_ _0291_ _0296_ _0297_ VGND
+ VGND VDPWR VDPWR _0332_ sky130_fd_sc_hd__a2111o_1
X_2103_ net164 _0750_ _0784_ _0794_ VGND VGND VDPWR VDPWR _0796_ sky130_fd_sc_hd__o211a_1
XFILLER_0_76_125 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[42\].gen_latches\[6\].p_latch net198 dig_ctrl_inst.latch_mem_inst.gclk\[42\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[42\]\[6\] sky130_fd_sc_hd__dlxtp_1
X_2034_ _0287_ _0719_ _0734_ _0738_ VGND VGND VDPWR VDPWR _0739_ sky130_fd_sc_hd__or4_4
X_1818_ dig_ctrl_inst.latch_mem_inst.RAM\[36\]\[4\] net96 net54 VGND VGND VDPWR VDPWR
+ _0526_ sky130_fd_sc_hd__and3_2
XFILLER_0_68_70 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
X_1749_ _0454_ _0455_ _0456_ _0457_ VGND VGND VDPWR VDPWR _0458_ sky130_fd_sc_hd__or4_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[31\].gen_latches\[4\].p_latch net208 dig_ctrl_inst.latch_mem_inst.gclk\[31\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[31\]\[4\] sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_68_573 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_169 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_331 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[20\].gen_latches\[2\].p_latch net228 dig_ctrl_inst.latch_mem_inst.gclk\[20\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[20\]\[2\] sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_51_473 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_29 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_6
Xdig_ctrl_inst.latch_mem_inst.gen_words\[58\].gen_latches\[0\].p_latch net246 dig_ctrl_inst.latch_mem_inst.gclk\[58\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[58\]\[0\] sky130_fd_sc_hd__dlxtp_1
X_1465_ dig_ctrl_inst.spi_addr\[3\] _0185_ _0191_ dig_ctrl_inst.spi_addr\[4\] VGND
+ VGND VDPWR VDPWR _0194_ sky130_fd_sc_hd__a31o_1
Xfanout119 _1129_ VGND VGND VDPWR VDPWR net119 sky130_fd_sc_hd__clkbuf_4
Xfanout108 _1134_ VGND VGND VDPWR VDPWR net108 sky130_fd_sc_hd__buf_4
X_1603_ dig_ctrl_inst.latch_mem_inst.RAM\[21\]\[0\] _0124_ _0155_ dig_ctrl_inst.latch_mem_inst.RAM\[58\]\[0\]
+ VGND VGND VDPWR VDPWR _0315_ sky130_fd_sc_hd__a22o_1
X_1534_ net167 net166 VGND VGND VDPWR VDPWR _0247_ sky130_fd_sc_hd__or2_1
XFILLER_0_1_155 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_65_554 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2017_ dig_ctrl_inst.latch_mem_inst.RAM\[25\]\[7\] _0128_ _0139_ dig_ctrl_inst.latch_mem_inst.RAM\[39\]\[7\]
+ _0721_ VGND VGND VDPWR VDPWR _0722_ sky130_fd_sc_hd__a221o_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[46\].gen_latches\[7\].p_latch net183 dig_ctrl_inst.latch_mem_inst.gclk\[46\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[46\]\[7\] sky130_fd_sc_hd__dlxtp_1
X_1396_ net149 _0153_ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.data_we\[55\]
+ sky130_fd_sc_hd__and2_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[2\].gen_latches\[2\].p_latch net225 dig_ctrl_inst.latch_mem_inst.gclk\[2\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[2\]\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_64_106 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_147 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_19_Left_97 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[35\].gen_latches\[5\].p_latch net200 dig_ctrl_inst.latch_mem_inst.gclk\[35\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[35\]\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_13_272 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_8
Xdig_ctrl_inst.latch_mem_inst.gen_words\[24\].gen_latches\[3\].p_latch net216 dig_ctrl_inst.latch_mem_inst.gclk\[24\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[24\]\[3\] sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[11\].clock_gate clknet_leaf_1_clk dig_ctrl_inst.latch_mem_inst.data_we\[11\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.gen_gclk\[11\]._gclk sky130_fd_sc_hd__dlclkp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[13\].gen_latches\[1\].p_latch net236 dig_ctrl_inst.latch_mem_inst.gclk\[13\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[13\]\[1\] sky130_fd_sc_hd__dlxtp_1
X_1250_ net182 net297 _1027_ dig_ctrl_inst.cpu_inst.ip\[5\] VGND VGND VDPWR VDPWR
+ _1098_ sky130_fd_sc_hd__o211a_1
X_1181_ net182 net292 _1027_ dig_ctrl_inst.cpu_inst.ip\[3\] VGND VGND VDPWR VDPWR
+ _1029_ sky130_fd_sc_hd__o211a_4
XTAP_TAPCELL_ROW_62_535 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_278 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_53 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
X_1448_ dig_ctrl_inst.spi_receiver_inst.spi_cnt\[0\] _0181_ dig_ctrl_inst.spi_receiver_inst.spi_cnt\[1\]
+ VGND VGND VDPWR VDPWR _0183_ sky130_fd_sc_hd__a21oi_1
X_2497_ clknet_leaf_8_clk dig_ctrl_inst.cpu_inst.stb_o net180 VGND VGND VDPWR VDPWR
+ dig_ctrl_inst.stb_d sky130_fd_sc_hd__dfrtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[6\].gen_latches\[3\].p_latch net220 dig_ctrl_inst.latch_mem_inst.gclk\[6\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[6\]\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_4_41 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_253 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
X_1517_ _0228_ _0229_ VGND VGND VDPWR VDPWR _0230_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_2_179 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1379_ net148 net72 net51 VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.data_we\[46\]
+ sky130_fd_sc_hd__and3_2
XFILLER_0_33_334 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[39\].gen_latches\[6\].p_latch net191 dig_ctrl_inst.latch_mem_inst.gclk\[39\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[39\]\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_60_153 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[28\].gen_latches\[4\].p_latch net209 dig_ctrl_inst.latch_mem_inst.gclk\[28\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[28\]\[4\] sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[17\].gen_latches\[2\].p_latch net230 dig_ctrl_inst.latch_mem_inst.gclk\[17\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[17\]\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_28_139 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_259 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_109 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
X_2420_ clknet_leaf_9_clk _0028_ net141 VGND VGND VDPWR VDPWR dig_ctrl_inst.cpu_inst.arg1\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout90 net92 VGND VGND VDPWR VDPWR net90 sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_23_Left_101 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
X_2351_ dig_ctrl_inst.cpu_inst.port_o\[6\] net34 _0987_ VGND VGND VDPWR VDPWR _0101_
+ sky130_fd_sc_hd__mux2_1
X_1302_ net124 net88 VGND VGND VDPWR VDPWR _1142_ sky130_fd_sc_hd__and2_2
X_2282_ _1022_ _0175_ _0756_ VGND VGND VDPWR VDPWR _0967_ sky130_fd_sc_hd__and3_4
X_1233_ net259 net255 dig_ctrl_inst.cpu_inst.r2\[1\] VGND VGND VDPWR VDPWR _1081_
+ sky130_fd_sc_hd__and3b_1
XFILLER_0_35_74 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_32_Left_110 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
X_1164_ _1011_ VGND VGND VDPWR VDPWR _1012_ sky130_fd_sc_hd__inv_2
X_1997_ dig_ctrl_inst.latch_mem_inst.RAM\[58\]\[7\] net85 net49 VGND VGND VDPWR VDPWR
+ _0702_ sky130_fd_sc_hd__and3_2
XFILLER_0_15_334 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_117 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[41\].clock_buffer dig_ctrl_inst.latch_mem_inst.gen_gclk\[41\]._gclk
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.gclk\[41\] sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_7_205 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_223 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_38_395 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_337 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_29_340 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1851_ dig_ctrl_inst.latch_mem_inst.RAM\[47\]\[4\] _0146_ _0152_ dig_ctrl_inst.latch_mem_inst.RAM\[54\]\[4\]
+ VGND VGND VDPWR VDPWR _0559_ sky130_fd_sc_hd__a22o_1
X_1920_ dig_ctrl_inst.latch_mem_inst.RAM\[43\]\[6\] net104 net91 net56 VGND VGND VDPWR
+ VDPWR _0626_ sky130_fd_sc_hd__and4_1
XFILLER_0_8_309 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_6
X_2403_ clknet_leaf_6_clk _0011_ net146 VGND VGND VDPWR VDPWR dig_ctrl_inst.cpu_inst.port_o\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_1782_ dig_ctrl_inst.latch_mem_inst.RAM\[19\]\[3\] net131 net103 net62 VGND VGND
+ VDPWR VDPWR _0491_ sky130_fd_sc_hd__and4_1
XFILLER_0_24_153 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_197 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_2334_ dig_ctrl_inst.spi_data_o\[6\] dig_ctrl_inst.spi_data_o\[7\] _0180_ VGND VGND
+ VDPWR VDPWR _0086_ sky130_fd_sc_hd__mux2_1
X_2196_ _0240_ _0884_ VGND VGND VDPWR VDPWR _0885_ sky130_fd_sc_hd__xnor2_1
X_2265_ _0236_ _0950_ VGND VGND VDPWR VDPWR _0951_ sky130_fd_sc_hd__xnor2_1
X_1216_ dig_ctrl_inst.cpu_inst.r3\[0\] net258 net254 VGND VGND VDPWR VDPWR _1064_
+ sky130_fd_sc_hd__and3_2
XTAP_TAPCELL_ROW_35_376 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_86 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_131 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_197 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
Xhold55 dig_ctrl_inst.spi_receiver_inst.synchronizer_spi_cs.pipe\[0\] VGND VGND VDPWR
+ VDPWR net337 sky130_fd_sc_hd__dlygate4sd3_1
Xhold66 dig_ctrl_inst.spi_data_i\[4\] VGND VGND VDPWR VDPWR net348 sky130_fd_sc_hd__dlygate4sd3_1
Xhold99 dig_ctrl_inst.cpu_inst.r2\[3\] VGND VGND VDPWR VDPWR net381 sky130_fd_sc_hd__dlygate4sd3_1
Xhold44 dig_ctrl_inst.latch_mem_inst.wdata\[5\] VGND VGND VDPWR VDPWR net326 sky130_fd_sc_hd__dlygate4sd3_1
Xhold77 dig_ctrl_inst.cpu_inst.r1\[4\] VGND VGND VDPWR VDPWR net359 sky130_fd_sc_hd__dlygate4sd3_1
Xhold88 dig_ctrl_inst.cpu_inst.r3\[3\] VGND VGND VDPWR VDPWR net370 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_26_321 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[61\].gen_latches\[4\].p_latch net210 dig_ctrl_inst.latch_mem_inst.gclk\[61\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[61\]\[4\] sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[50\].gen_latches\[2\].p_latch net228 dig_ctrl_inst.latch_mem_inst.gclk\[50\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[50\]\[2\] sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_7_Left_85 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_39 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XANTENNA_8 _0674_ VGND VGND VDPWR VDPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_457 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2050_ dig_ctrl_inst.cpu_inst.instr\[5\] _1012_ _1013_ net296 VGND VGND VDPWR VDPWR
+ _0743_ sky130_fd_sc_hd__o211a_2
XFILLER_0_29_223 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_1834_ dig_ctrl_inst.latch_mem_inst.RAM\[8\]\[4\] _1142_ _0539_ _0540_ _0541_ VGND
+ VGND VDPWR VDPWR _0542_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_32_357 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1903_ dig_ctrl_inst.latch_mem_inst.RAM\[18\]\[5\] net109 net61 VGND VGND VDPWR VDPWR
+ _0610_ sky130_fd_sc_hd__and3_2
X_1765_ dig_ctrl_inst.latch_mem_inst.RAM\[24\]\[3\] net86 net67 VGND VGND VDPWR VDPWR
+ _0474_ sky130_fd_sc_hd__and3_2
X_1696_ dig_ctrl_inst.latch_mem_inst.RAM\[27\]\[2\] net105 net91 net66 VGND VGND VDPWR
+ VDPWR _0406_ sky130_fd_sc_hd__and4_1
X_2317_ dig_ctrl_inst.spi_receiver_inst.spi_cs_sync dig_ctrl_inst.spi_receiver_inst.spi_sclk_delayed
+ dig_ctrl_inst.spi_receiver_inst.spi_sclk_sync VGND VGND VDPWR VDPWR _0978_ sky130_fd_sc_hd__or3b_1
XFILLER_0_32_3 VDPWR VGND VDPWR VGND sky130_ef_sc_hd__decap_12
X_2248_ _0933_ _0934_ VGND VGND VDPWR VDPWR _0935_ sky130_fd_sc_hd__nand2_1
X_2179_ _0867_ _0868_ VGND VGND VDPWR VDPWR _0869_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_23_302 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput34 net34 VGND VGND VDPWR VDPWR uo_out[6] sky130_fd_sc_hd__buf_2
Xoutput23 net23 VGND VGND VDPWR VDPWR port_ms_o[6] sky130_fd_sc_hd__buf_2
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[16\].clock_gate clknet_leaf_15_clk dig_ctrl_inst.latch_mem_inst.data_we\[16\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.gen_gclk\[16\]._gclk sky130_fd_sc_hd__dlclkp_1
XTAP_TAPCELL_ROW_46_438 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[54\].gen_latches\[3\].p_latch net216 dig_ctrl_inst.latch_mem_inst.gclk\[54\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[54\]\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_5_109 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
X_1481_ dig_ctrl_inst.stb_d dig_ctrl_inst.stb_dd _1039_ VGND VGND VDPWR VDPWR _0200_
+ sky130_fd_sc_hd__mux2_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[43\].gen_latches\[1\].p_latch net234 dig_ctrl_inst.latch_mem_inst.gclk\[43\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[43\]\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_1_337 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
X_1550_ net161 net163 VGND VGND VDPWR VDPWR _0263_ sky130_fd_sc_hd__and2b_1
X_2033_ _0737_ _0735_ _0736_ _0720_ VGND VGND VDPWR VDPWR _0738_ sky130_fd_sc_hd__or4_4
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[34\].clock_buffer dig_ctrl_inst.latch_mem_inst.gen_gclk\[34\]._gclk
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.gclk\[34\] sky130_fd_sc_hd__clkbuf_4
X_2102_ dig_ctrl_inst.cpu_inst.data\[0\] _0743_ _0747_ net164 VGND VGND VDPWR VDPWR
+ _0795_ sky130_fd_sc_hd__a22oi_1
X_1748_ dig_ctrl_inst.latch_mem_inst.RAM\[18\]\[3\] _0121_ _0136_ dig_ctrl_inst.latch_mem_inst.RAM\[34\]\[3\]
+ VGND VGND VDPWR VDPWR _0457_ sky130_fd_sc_hd__a22o_1
XFILLER_0_25_281 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_63 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
X_1817_ dig_ctrl_inst.latch_mem_inst.RAM\[10\]\[4\] net121 net84 VGND VGND VDPWR VDPWR
+ _0525_ sky130_fd_sc_hd__and3_2
XFILLER_0_68_93 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_1679_ dig_ctrl_inst.latch_mem_inst.RAM\[13\]\[1\] _0114_ _0342_ _0343_ _0364_ VGND
+ VGND VDPWR VDPWR _0390_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_68_574 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[20\].gen_latches\[6\].p_latch net198 dig_ctrl_inst.latch_mem_inst.gclk\[20\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[20\]\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_64_29 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_8
Xdig_ctrl_inst.latch_mem_inst.gen_words\[58\].gen_latches\[4\].p_latch net212 dig_ctrl_inst.latch_mem_inst.gclk\[58\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[58\]\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_13_55 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_1602_ dig_ctrl_inst.latch_mem_inst.RAM\[50\]\[0\] net112 net50 _0129_ dig_ctrl_inst.latch_mem_inst.RAM\[26\]\[0\]
+ VGND VGND VDPWR VDPWR _0314_ sky130_fd_sc_hd__a32o_1
XFILLER_0_22_251 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[47\].gen_latches\[2\].p_latch net225 dig_ctrl_inst.latch_mem_inst.gclk\[47\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[47\]\[2\] sky130_fd_sc_hd__dlxtp_1
X_1464_ _0193_ _0192_ dig_ctrl_inst.spi_addr\[3\] VGND VGND VDPWR VDPWR _0008_ sky130_fd_sc_hd__mux2_1
X_1533_ net167 net166 VGND VGND VDPWR VDPWR _0246_ sky130_fd_sc_hd__nand2_1
X_1395_ net102 net99 net42 VGND VGND VDPWR VDPWR _0153_ sky130_fd_sc_hd__and3_4
Xfanout109 net112 VGND VGND VDPWR VDPWR net109 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_65_555 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_51 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_8
X_2016_ dig_ctrl_inst.latch_mem_inst.RAM\[27\]\[7\] _0130_ _0152_ dig_ctrl_inst.latch_mem_inst.RAM\[54\]\[7\]
+ VGND VGND VDPWR VDPWR _0721_ sky130_fd_sc_hd__a22o_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[36\].gen_latches\[0\].p_latch net246 dig_ctrl_inst.latch_mem_inst.gclk\[36\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[36\]\[0\] sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[2\].gen_latches\[6\].p_latch net193 dig_ctrl_inst.latch_mem_inst.gclk\[2\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[2\]\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_60_313 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_223 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_500 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[24\].gen_latches\[7\].p_latch net185 dig_ctrl_inst.latch_mem_inst.gclk\[24\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[24\]\[7\] sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[13\].gen_latches\[5\].p_latch net201 dig_ctrl_inst.latch_mem_inst.gclk\[13\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[13\]\[5\] sky130_fd_sc_hd__dlxtp_1
X_1180_ net297 net182 _1027_ VGND VGND VDPWR VDPWR _1028_ sky130_fd_sc_hd__o21a_1
XPHY_EDGE_ROW_20_Left_98 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_19_279 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_536 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_12_clk clknet_1_0__leaf_clk VGND VGND VDPWR VDPWR clknet_leaf_12_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_10_221 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
X_1516_ _0167_ net138 VGND VGND VDPWR VDPWR _0229_ sky130_fd_sc_hd__nor2_1
X_1447_ dig_ctrl_inst.spi_receiver_inst.spi_cnt\[0\] dig_ctrl_inst.spi_receiver_inst.spi_cnt\[1\]
+ _0181_ VGND VGND VDPWR VDPWR _0182_ sky130_fd_sc_hd__and3_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[6\].gen_latches\[7\].p_latch net187 dig_ctrl_inst.latch_mem_inst.gclk\[6\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[6\]\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_49_95 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
X_2496_ clknet_leaf_7_clk net343 net180 VGND VGND VDPWR VDPWR dig_ctrl_inst.stb_dd
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_287 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_298 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
X_1378_ net149 _0145_ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.data_we\[45\]
+ sky130_fd_sc_hd__and2_1
Xfanout91 net92 VGND VGND VDPWR VDPWR net91 sky130_fd_sc_hd__clkbuf_2
Xfanout80 net81 VGND VGND VDPWR VDPWR net80 sky130_fd_sc_hd__buf_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[17\].gen_latches\[6\].p_latch net195 dig_ctrl_inst.latch_mem_inst.gclk\[17\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[17\]\[6\] sky130_fd_sc_hd__dlxtp_1
X_2350_ dig_ctrl_inst.cpu_inst.port_o\[5\] net33 _0987_ VGND VGND VDPWR VDPWR _0100_
+ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_1_clk clknet_1_1__leaf_clk VGND VGND VDPWR VDPWR clknet_leaf_1_clk sky130_fd_sc_hd__clkbuf_8
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[27\].clock_buffer dig_ctrl_inst.latch_mem_inst.gen_gclk\[27\]._gclk
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.gclk\[27\] sky130_fd_sc_hd__clkbuf_4
X_1301_ net305 _1078_ _1093_ _1062_ _1048_ VGND VGND VDPWR VDPWR _1141_ sky130_fd_sc_hd__a2111oi_2
X_2281_ _0963_ _0966_ _0949_ VGND VGND VDPWR VDPWR _0052_ sky130_fd_sc_hd__a21oi_1
X_1232_ net258 net255 dig_ctrl_inst.cpu_inst.r3\[1\] VGND VGND VDPWR VDPWR _1080_
+ sky130_fd_sc_hd__and3_2
XFILLER_0_35_97 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_1163_ net258 net254 VGND VGND VDPWR VDPWR _1011_ sky130_fd_sc_hd__nand2b_2
XFILLER_0_51_96 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
X_1996_ dig_ctrl_inst.latch_mem_inst.RAM\[47\]\[7\] _0146_ _0148_ dig_ctrl_inst.latch_mem_inst.RAM\[49\]\[7\]
+ VGND VGND VDPWR VDPWR _0701_ sky130_fd_sc_hd__a22o_1
XFILLER_0_62_3 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_251 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_240 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_7_206 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2479_ clknet_leaf_2_clk _0085_ net180 VGND VGND VDPWR VDPWR dig_ctrl_inst.spi_data_o\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_65_279 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_202 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
Xclkload0 clknet_1_0__leaf_clk VGND VGND VDPWR VDPWR clkload0/Y sky130_fd_sc_hd__inv_8
XTAP_TAPCELL_ROW_29_341 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[23\].clock_gate clknet_leaf_12_clk dig_ctrl_inst.latch_mem_inst.data_we\[23\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.gen_gclk\[23\]._gclk sky130_fd_sc_hd__dlclkp_1
X_1850_ _0555_ _0556_ _0557_ VGND VGND VDPWR VDPWR _0558_ sky130_fd_sc_hd__or3_1
XFILLER_0_21_44 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
X_1781_ dig_ctrl_inst.latch_mem_inst.RAM\[16\]\[3\] _0119_ _0487_ _0488_ _0489_ VGND
+ VGND VDPWR VDPWR _0490_ sky130_fd_sc_hd__a2111o_1
X_2402_ clknet_leaf_6_clk _0000_ net145 VGND VGND VDPWR VDPWR dig_ctrl_inst.cpu_inst.port_stb_o
+ sky130_fd_sc_hd__dfrtp_4
X_2333_ dig_ctrl_inst.spi_data_o\[5\] dig_ctrl_inst.spi_data_o\[6\] _0180_ VGND VGND
+ VDPWR VDPWR _0085_ sky130_fd_sc_hd__mux2_1
X_1215_ _1047_ net135 VGND VGND VDPWR VDPWR _1063_ sky130_fd_sc_hd__nor2_1
X_2195_ _0252_ _0864_ _0249_ VGND VGND VDPWR VDPWR _0884_ sky130_fd_sc_hd__o21a_1
X_2264_ _0230_ _0927_ _0228_ VGND VGND VDPWR VDPWR _0950_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_62_51 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_279 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_35_377 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_321 VDPWR VGND VDPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_290 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
X_1979_ dig_ctrl_inst.latch_mem_inst.RAM\[0\]\[6\] _0288_ _0671_ _0684_ VGND VGND
+ VDPWR VDPWR _0685_ sky130_fd_sc_hd__o22a_4
Xhold56 dig_ctrl_inst.synchronizer_port_i_inst\[6\].pipe\[0\] VGND VGND VDPWR VDPWR
+ net338 sky130_fd_sc_hd__dlygate4sd3_1
Xhold45 dig_ctrl_inst.latch_mem_inst.wdata\[1\] VGND VGND VDPWR VDPWR net327 sky130_fd_sc_hd__dlygate4sd3_1
Xhold89 dig_ctrl_inst.cpu_inst.r2\[2\] VGND VGND VDPWR VDPWR net371 sky130_fd_sc_hd__dlygate4sd3_1
Xhold67 dig_ctrl_inst.cpu_inst.prev_state\[1\] VGND VGND VDPWR VDPWR net349 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_26_322 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold78 dig_ctrl_inst.cpu_inst.r3\[0\] VGND VGND VDPWR VDPWR net360 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_51_Left_129 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XANTENNA_9 _1136_ VGND VGND VDPWR VDPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_60_Left_138 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[50\].gen_latches\[6\].p_latch net192 dig_ctrl_inst.latch_mem_inst.gclk\[50\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[50\]\[6\] sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_49_458 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1902_ dig_ctrl_inst.latch_mem_inst.RAM\[49\]\[5\] net131 net114 net42 VGND VGND
+ VDPWR VDPWR _0609_ sky130_fd_sc_hd__and4_1
X_1764_ dig_ctrl_inst.latch_mem_inst.RAM\[11\]\[3\] _1145_ _0470_ _0471_ _0472_ VGND
+ VGND VDPWR VDPWR _0473_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_32_358 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1833_ dig_ctrl_inst.latch_mem_inst.RAM\[28\]\[4\] net77 net65 VGND VGND VDPWR VDPWR
+ _0541_ sky130_fd_sc_hd__and3_2
X_1695_ dig_ctrl_inst.latch_mem_inst.RAM\[19\]\[2\] net132 net107 net69 VGND VGND
+ VDPWR VDPWR _0405_ sky130_fd_sc_hd__and4_1
X_2316_ net364 _0975_ _0977_ VGND VGND VDPWR VDPWR _0076_ sky130_fd_sc_hd__mux2_1
X_2247_ net138 _0911_ VGND VGND VDPWR VDPWR _0934_ sky130_fd_sc_hd__nand2_1
X_2178_ net169 _0842_ VGND VGND VDPWR VDPWR _0868_ sky130_fd_sc_hd__nand2_1
XFILLER_0_25_3 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_23_303 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput35 net35 VGND VGND VDPWR VDPWR uo_out[7] sky130_fd_sc_hd__buf_2
Xoutput24 net24 VGND VGND VDPWR VDPWR port_ms_o[7] sky130_fd_sc_hd__buf_2
XFILLER_0_50_208 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_190 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_46_439 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_19_Right_19 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[54\].gen_latches\[7\].p_latch net189 dig_ctrl_inst.latch_mem_inst.gclk\[54\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[54\]\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_1_305 VDPWR VGND VDPWR VGND sky130_ef_sc_hd__decap_12
X_1480_ _1023_ _0175_ _0198_ VGND VGND VDPWR VDPWR _0199_ sky130_fd_sc_hd__and3_2
XPHY_EDGE_ROW_28_Right_28 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_31 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_37_Right_37 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[43\].gen_latches\[5\].p_latch net202 dig_ctrl_inst.latch_mem_inst.gclk\[43\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[43\]\[5\] sky130_fd_sc_hd__dlxtp_1
X_2032_ dig_ctrl_inst.latch_mem_inst.RAM\[55\]\[7\] _0153_ _0687_ _0695_ _0706_ VGND
+ VGND VDPWR VDPWR _0737_ sky130_fd_sc_hd__a2111o_1
X_2101_ _0786_ _0791_ net158 VGND VGND VDPWR VDPWR _0794_ sky130_fd_sc_hd__mux2_1
XFILLER_0_57_341 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_64 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[32\].gen_latches\[3\].p_latch net217 dig_ctrl_inst.latch_mem_inst.gclk\[32\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[32\]\[3\] sky130_fd_sc_hd__dlxtp_1
X_1747_ dig_ctrl_inst.latch_mem_inst.RAM\[30\]\[3\] net73 net70 _0156_ dig_ctrl_inst.latch_mem_inst.RAM\[59\]\[3\]
+ VGND VGND VDPWR VDPWR _0456_ sky130_fd_sc_hd__a32o_1
XPHY_EDGE_ROW_46_Right_46 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_263 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
X_1678_ dig_ctrl_inst.latch_mem_inst.RAM\[31\]\[1\] _0132_ _0345_ _0346_ _0354_ VGND
+ VGND VDPWR VDPWR _0389_ sky130_fd_sc_hd__a2111o_1
X_1816_ dig_ctrl_inst.latch_mem_inst.RAM\[19\]\[4\] net133 net104 net64 VGND VGND
+ VDPWR VDPWR _0524_ sky130_fd_sc_hd__and4_1
XPHY_EDGE_ROW_55_Right_55 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[21\].gen_latches\[1\].p_latch net233 dig_ctrl_inst.latch_mem_inst.gclk\[21\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[21\]\[1\] sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_68_575 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_64_Right_64 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_271 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_73_Right_73 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_59_520 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[2\].clock_gate clknet_leaf_12_clk dig_ctrl_inst.latch_mem_inst.data_we\[2\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.gen_gclk\[2\]._gclk sky130_fd_sc_hd__dlclkp_1
XFILLER_0_58_127 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_341 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_1601_ dig_ctrl_inst.latch_mem_inst.RAM\[31\]\[0\] _0132_ _0277_ dig_ctrl_inst.latch_mem_inst.RAM\[4\]\[0\]
+ _0312_ VGND VGND VDPWR VDPWR _0313_ sky130_fd_sc_hd__a221o_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[3\].gen_latches\[1\].p_latch net238 dig_ctrl_inst.latch_mem_inst.gclk\[3\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[3\]\[1\] sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[47\].gen_latches\[6\].p_latch net197 dig_ctrl_inst.latch_mem_inst.gclk\[47\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[47\]\[6\] sky130_fd_sc_hd__dlxtp_1
X_1532_ _0244_ _0237_ _0240_ VGND VGND VDPWR VDPWR _0245_ sky130_fd_sc_hd__or3b_1
X_1463_ _0186_ _0191_ VGND VGND VDPWR VDPWR _0193_ sky130_fd_sc_hd__and2_1
XFILLER_0_38_97 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
X_1394_ net148 net93 net42 VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.data_we\[54\]
+ sky130_fd_sc_hd__and3_2
XTAP_TAPCELL_ROW_65_556 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2015_ _0692_ _0693_ _0694_ _0705_ VGND VGND VDPWR VDPWR _0720_ sky130_fd_sc_hd__or4_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[36\].gen_latches\[4\].p_latch net208 dig_ctrl_inst.latch_mem_inst.gclk\[36\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[36\]\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_72_141 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_279 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[25\].gen_latches\[2\].p_latch net224 dig_ctrl_inst.latch_mem_inst.gclk\[25\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[25\]\[2\] sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_56_501 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdig_ctrl_inst.latch_mem_inst.gen_input_latches\[2\].n_latch dig_ctrl_inst.data_out\[2\]
+ clknet_leaf_8_clk VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.wdata\[2\]
+ sky130_fd_sc_hd__dlxtn_1
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[28\].clock_gate clknet_leaf_0_clk dig_ctrl_inst.latch_mem_inst.data_we\[28\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.gen_gclk\[28\]._gclk sky130_fd_sc_hd__dlclkp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[14\].gen_latches\[0\].p_latch net247 dig_ctrl_inst.latch_mem_inst.gclk\[14\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[14\]\[0\] sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_62_537 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[7\].gen_latches\[2\].p_latch net229 dig_ctrl_inst.latch_mem_inst.gclk\[7\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[7\]\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_54_141 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_130 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_193 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_77 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[30\].clock_gate clknet_leaf_0_clk dig_ctrl_inst.latch_mem_inst.data_we\[30\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.gen_gclk\[30\]._gclk sky130_fd_sc_hd__dlclkp_1
X_2495_ clknet_leaf_5_clk _0094_ net179 VGND VGND VDPWR VDPWR dig_ctrl_inst.spi_data_i\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_64_7 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_1515_ _0167_ net138 VGND VGND VDPWR VDPWR _0228_ sky130_fd_sc_hd__and2_1
X_1446_ dig_ctrl_inst.spi_receiver_inst.spi_cnt\[0\] _0180_ VGND VGND VDPWR VDPWR
+ _0002_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_65_51 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
X_1377_ net115 net80 net52 VGND VGND VDPWR VDPWR _0145_ sky130_fd_sc_hd__and3_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[29\].gen_latches\[3\].p_latch net221 dig_ctrl_inst.latch_mem_inst.gclk\[29\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[29\]\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_5_271 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_76_618 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[18\].gen_latches\[1\].p_latch net232 dig_ctrl_inst.latch_mem_inst.gclk\[18\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[18\]\[1\] sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_1_170 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout70 net71 VGND VGND VDPWR VDPWR net70 sky130_fd_sc_hd__buf_2
Xfanout92 _1140_ VGND VGND VDPWR VDPWR net92 sky130_fd_sc_hd__buf_4
XFILLER_0_36_141 VDPWR VGND VDPWR VGND sky130_ef_sc_hd__decap_12
Xfanout81 _1146_ VGND VGND VDPWR VDPWR net81 sky130_fd_sc_hd__buf_2
XFILLER_0_51_155 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_1300_ net136 net135 VGND VGND VDPWR VDPWR _1140_ sky130_fd_sc_hd__nor2_1
X_1162_ net248 dig_ctrl_inst.cpu_inst.cpu_state\[2\] dig_ctrl_inst.cpu_inst.cpu_state\[1\]
+ VGND VGND VDPWR VDPWR _1010_ sky130_fd_sc_hd__nor3b_2
X_1231_ _1026_ net182 _1027_ dig_ctrl_inst.cpu_inst.ip\[1\] VGND VGND VDPWR VDPWR
+ _1079_ sky130_fd_sc_hd__o211a_1
X_2280_ _0754_ _0964_ _0965_ _0756_ net41 VGND VGND VDPWR VDPWR _0966_ sky130_fd_sc_hd__o221a_1
XFILLER_0_35_21 VDPWR VGND VDPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_44 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_99 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_188 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_122 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_111 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
X_1995_ dig_ctrl_inst.latch_mem_inst.RAM\[36\]\[7\] net96 net54 VGND VGND VDPWR VDPWR
+ _0700_ sky130_fd_sc_hd__and3_2
X_2478_ clknet_leaf_4_clk _0084_ net172 VGND VGND VDPWR VDPWR dig_ctrl_inst.spi_data_o\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_55_3 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_7_207 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1429_ net255 dig_ctrl_inst.cpu_inst.r1\[7\] VGND VGND VDPWR VDPWR _0170_ sky130_fd_sc_hd__and2b_1
XFILLER_0_65_225 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
Xclkload1 clknet_leaf_10_clk VGND VGND VDPWR VDPWR clkload1/Y sky130_fd_sc_hd__inv_16
XFILLER_0_18_141 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_317 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
Xfanout260 net261 VGND VGND VDPWR VDPWR net260 sky130_fd_sc_hd__buf_4
XFILLER_0_71_228 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_1780_ dig_ctrl_inst.latch_mem_inst.RAM\[10\]\[3\] net121 net294 VGND VGND VDPWR
+ VDPWR _0489_ sky130_fd_sc_hd__and3_2
X_2401_ clknet_leaf_4_clk _0010_ net176 VGND VGND VDPWR VDPWR dig_ctrl_inst.spi_addr\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_2332_ dig_ctrl_inst.spi_data_o\[4\] dig_ctrl_inst.spi_data_o\[5\] _0180_ VGND VGND
+ VDPWR VDPWR _0084_ sky130_fd_sc_hd__mux2_1
XFILLER_0_41_9 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_2194_ dig_ctrl_inst.cpu_inst.r0\[4\] _0758_ VGND VGND VDPWR VDPWR _0883_ sky130_fd_sc_hd__nor2_1
X_1214_ _1049_ _1055_ _1061_ dig_ctrl_inst.spi_addr\[2\] _1002_ VGND VGND VDPWR VDPWR
+ _1062_ sky130_fd_sc_hd__o32a_4
XFILLER_0_46_97 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
X_2263_ dig_ctrl_inst.cpu_inst.r0\[7\] net41 VGND VGND VDPWR VDPWR _0949_ sky130_fd_sc_hd__nor2_1
XFILLER_0_1_55 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_206 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_85 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_333 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[62\].gen_latches\[3\].p_latch net221 dig_ctrl_inst.latch_mem_inst.gclk\[62\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[62\]\[3\] sky130_fd_sc_hd__dlxtp_1
X_1978_ _0287_ _0674_ _0679_ _0683_ VGND VGND VDPWR VDPWR _0684_ sky130_fd_sc_hd__or4_4
Xhold57 dig_ctrl_inst.synchronizer_port_i_inst\[7\].pipe\[0\] VGND VGND VDPWR VDPWR
+ net339 sky130_fd_sc_hd__dlygate4sd3_1
Xhold68 dig_ctrl_inst.spi_data_i\[6\] VGND VGND VDPWR VDPWR net350 sky130_fd_sc_hd__dlygate4sd3_1
Xhold46 dig_ctrl_inst.latch_mem_inst.wdata\[7\] VGND VGND VDPWR VDPWR net328 sky130_fd_sc_hd__dlygate4sd3_1
Xhold79 dig_ctrl_inst.cpu_inst.r1\[6\] VGND VGND VDPWR VDPWR net361 sky130_fd_sc_hd__dlygate4sd3_1
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[7\].clock_gate clknet_leaf_1_clk dig_ctrl_inst.latch_mem_inst.data_we\[7\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.gen_gclk\[7\]._gclk sky130_fd_sc_hd__dlclkp_1
XTAP_TAPCELL_ROW_26_323 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[51\].gen_latches\[1\].p_latch net233 dig_ctrl_inst.latch_mem_inst.gclk\[51\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[51\]\[1\] sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_49_459 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1832_ dig_ctrl_inst.latch_mem_inst.RAM\[52\]\[4\] net96 net45 VGND VGND VDPWR VDPWR
+ _0540_ sky130_fd_sc_hd__and3_2
XTAP_TAPCELL_ROW_32_359 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_236 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_225 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
X_1901_ dig_ctrl_inst.latch_mem_inst.RAM\[41\]\[5\] net114 net90 net52 VGND VGND VDPWR
+ VDPWR _0608_ sky130_fd_sc_hd__and4_1
X_1763_ dig_ctrl_inst.latch_mem_inst.RAM\[51\]\[3\] net132 net106 net49 VGND VGND
+ VDPWR VDPWR _0472_ sky130_fd_sc_hd__and4_1
XFILLER_0_52_250 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
X_1694_ dig_ctrl_inst.latch_mem_inst.RAM\[43\]\[2\] _0143_ VGND VGND VDPWR VDPWR _0404_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_57_52 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
X_2315_ net352 _0974_ _0977_ VGND VGND VDPWR VDPWR _0075_ sky130_fd_sc_hd__mux2_1
X_2246_ net138 _0911_ VGND VGND VDPWR VDPWR _0933_ sky130_fd_sc_hd__or2_1
X_2177_ net169 _0842_ VGND VGND VDPWR VDPWR _0867_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_23_304 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput25 net25 VGND VGND VDPWR VDPWR uio_out[2] sky130_fd_sc_hd__buf_2
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[59\].clock_buffer dig_ctrl_inst.latch_mem_inst.gen_gclk\[59\]._gclk
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.gclk\[59\] sky130_fd_sc_hd__clkbuf_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[55\].gen_latches\[2\].p_latch net224 dig_ctrl_inst.latch_mem_inst.gclk\[55\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[55\]\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_58_309 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[44\].gen_latches\[0\].p_latch net244 dig_ctrl_inst.latch_mem_inst.gclk\[44\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[44\]\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_34_250 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_317 VDPWR VGND VDPWR VGND sky130_ef_sc_hd__decap_12
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[35\].clock_gate clknet_leaf_16_clk dig_ctrl_inst.latch_mem_inst.data_we\[35\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.gen_gclk\[35\]._gclk sky130_fd_sc_hd__dlclkp_1
X_2100_ _1016_ _0745_ VGND VGND VDPWR VDPWR _0793_ sky130_fd_sc_hd__or2_2
X_2031_ _1145_ dig_ctrl_inst.latch_mem_inst.RAM\[11\]\[7\] _0691_ _0698_ _0703_ VGND
+ VGND VDPWR VDPWR _0736_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_27_55 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_209 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
X_1815_ dig_ctrl_inst.latch_mem_inst.RAM\[31\]\[4\] _0132_ _0520_ _0521_ _0522_ VGND
+ VGND VDPWR VDPWR _0523_ sky130_fd_sc_hd__a2111o_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[32\].gen_latches\[7\].p_latch net187 dig_ctrl_inst.latch_mem_inst.gclk\[32\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[32\]\[7\] sky130_fd_sc_hd__dlxtp_1
X_1746_ dig_ctrl_inst.latch_mem_inst.RAM\[22\]\[3\] _0125_ _0159_ dig_ctrl_inst.latch_mem_inst.RAM\[62\]\[3\]
+ VGND VGND VDPWR VDPWR _0455_ sky130_fd_sc_hd__a22o_1
XFILLER_0_40_253 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_1677_ dig_ctrl_inst.latch_mem_inst.RAM\[15\]\[1\] _0117_ _0143_ dig_ctrl_inst.latch_mem_inst.RAM\[43\]\[1\]
+ _0367_ VGND VGND VDPWR VDPWR _0388_ sky130_fd_sc_hd__a221o_1
XFILLER_0_4_166 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_2229_ _0241_ _0243_ _0787_ _0914_ _0916_ VGND VGND VDPWR VDPWR _0917_ sky130_fd_sc_hd__o311a_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[21\].gen_latches\[5\].p_latch net202 dig_ctrl_inst.latch_mem_inst.gclk\[21\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[21\]\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_75_183 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[59\].gen_latches\[3\].p_latch net222 dig_ctrl_inst.latch_mem_inst.gclk\[59\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[59\]\[3\] sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_59_521 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_3 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[10\].gen_latches\[3\].p_latch net217 dig_ctrl_inst.latch_mem_inst.gclk\[10\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[10\]\[3\] sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[48\].gen_latches\[1\].p_latch net236 dig_ctrl_inst.latch_mem_inst.gclk\[48\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[48\]\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_66_183 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_301 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_1462_ _0190_ _0192_ VGND VGND VDPWR VDPWR _0007_ sky130_fd_sc_hd__and2_1
X_1600_ dig_ctrl_inst.latch_mem_inst.RAM\[30\]\[0\] net74 net69 _0142_ dig_ctrl_inst.latch_mem_inst.RAM\[42\]\[0\]
+ VGND VGND VDPWR VDPWR _0312_ sky130_fd_sc_hd__a32o_1
XFILLER_0_1_169 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_1531_ _0241_ _0243_ VGND VGND VDPWR VDPWR _0244_ sky130_fd_sc_hd__nor2_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[3\].gen_latches\[5\].p_latch net201 dig_ctrl_inst.latch_mem_inst.gclk\[3\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[3\]\[5\] sky130_fd_sc_hd__dlxtp_1
X_1393_ net94 net46 VGND VGND VDPWR VDPWR _0152_ sky130_fd_sc_hd__and2_2
X_2014_ dig_ctrl_inst.latch_mem_inst.RAM\[8\]\[7\] _1142_ _0142_ dig_ctrl_inst.latch_mem_inst.RAM\[42\]\[7\]
+ _0718_ VGND VGND VDPWR VDPWR _0719_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_65_557 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_97 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_139 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_117 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
Xhold110 net18 VGND VGND VDPWR VDPWR net392 sky130_fd_sc_hd__dlygate4sd3_1
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[30\].clock_buffer dig_ctrl_inst.latch_mem_inst.gen_gclk\[30\]._gclk
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.gclk\[30\] sky130_fd_sc_hd__clkbuf_4
X_1729_ _0432_ _0436_ _0437_ _0438_ VGND VGND VDPWR VDPWR _0439_ sky130_fd_sc_hd__or4_1
XFILLER_0_13_297 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_56_502 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdig_ctrl_inst.latch_mem_inst.gen_input_latches\[6\].n_latch dig_ctrl_inst.data_out\[6\]
+ clknet_leaf_8_clk VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.wdata\[6\]
+ sky130_fd_sc_hd__dlxtn_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[25\].gen_latches\[6\].p_latch net194 dig_ctrl_inst.latch_mem_inst.gclk\[25\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[25\]\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_48_161 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[14\].gen_latches\[4\].p_latch net213 dig_ctrl_inst.latch_mem_inst.gclk\[14\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[14\]\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_51_337 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_62_538 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_190 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_23 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_89 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_70_582 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_153 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_217 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[7\].gen_latches\[6\].p_latch net198 dig_ctrl_inst.latch_mem_inst.gclk\[7\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[7\]\[6\] sky130_fd_sc_hd__dlxtp_1
X_2494_ clknet_leaf_6_clk _0093_ net179 VGND VGND VDPWR VDPWR dig_ctrl_inst.spi_data_i\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_1445_ _0180_ VGND VGND VDPWR VDPWR _0181_ sky130_fd_sc_hd__inv_2
X_1514_ net265 net262 dig_ctrl_inst.cpu_inst.r0\[6\] _0225_ _0226_ VGND VGND VDPWR
+ VDPWR _0227_ sky130_fd_sc_hd__o32a_1
XFILLER_0_4_11 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_63 VDPWR VGND VDPWR VGND sky130_ef_sc_hd__decap_12
X_1376_ net156 net78 net58 VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.data_we\[44\]
+ sky130_fd_sc_hd__and3_2
XTAP_TAPCELL_ROW_18_270 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[29\].gen_latches\[7\].p_latch net187 dig_ctrl_inst.latch_mem_inst.gclk\[29\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[29\]\[7\] sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_76_619 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_109 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_1_171 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[18\].gen_latches\[5\].p_latch net199 dig_ctrl_inst.latch_mem_inst.gclk\[18\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[18\]\[5\] sky130_fd_sc_hd__dlxtp_1
Xfanout82 _1146_ VGND VGND VDPWR VDPWR net82 sky130_fd_sc_hd__clkbuf_4
Xfanout60 _0133_ VGND VGND VDPWR VDPWR net60 sky130_fd_sc_hd__buf_6
Xfanout71 _0118_ VGND VGND VDPWR VDPWR net71 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_36_153 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
Xfanout93 net95 VGND VGND VDPWR VDPWR net93 sky130_fd_sc_hd__buf_2
X_1230_ dig_ctrl_inst.spi_addr\[0\] _1002_ VGND VGND VDPWR VDPWR _1078_ sky130_fd_sc_hd__or2_2
X_1161_ dig_ctrl_inst.cpu_inst.cpu_state\[1\] dig_ctrl_inst.cpu_inst.cpu_state\[2\]
+ net248 VGND VGND VDPWR VDPWR _1009_ sky130_fd_sc_hd__nor3b_1
XFILLER_0_35_55 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_1994_ dig_ctrl_inst.latch_mem_inst.RAM\[46\]\[7\] net75 net55 VGND VGND VDPWR VDPWR
+ _0699_ sky130_fd_sc_hd__and3_2
XFILLER_0_42_145 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_307 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_253 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_337 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
X_2477_ clknet_leaf_4_clk _0083_ net172 VGND VGND VDPWR VDPWR dig_ctrl_inst.spi_data_o\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_48_3 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_7_208 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1428_ net258 net254 dig_ctrl_inst.cpu_inst.r2\[7\] VGND VGND VDPWR VDPWR _0169_
+ sky130_fd_sc_hd__and3b_1
X_1359_ net131 net102 net51 VGND VGND VDPWR VDPWR _0137_ sky130_fd_sc_hd__and3_4
Xclkload2 clknet_leaf_11_clk VGND VGND VDPWR VDPWR clkload2/Y sky130_fd_sc_hd__inv_12
XFILLER_0_18_197 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
Xfanout250 net251 VGND VGND VDPWR VDPWR net250 sky130_fd_sc_hd__clkbuf_2
Xfanout261 dig_ctrl_inst.cpu_inst.arg1\[0\] VGND VGND VDPWR VDPWR net261 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_56_215 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_2400_ clknet_leaf_4_clk _0009_ net176 VGND VGND VDPWR VDPWR dig_ctrl_inst.spi_addr\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_35 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_57 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_6
X_2331_ dig_ctrl_inst.spi_data_o\[3\] dig_ctrl_inst.spi_data_o\[4\] _0180_ VGND VGND
+ VDPWR VDPWR _0083_ sky130_fd_sc_hd__mux2_1
X_1213_ _1039_ _1060_ net249 VGND VGND VDPWR VDPWR _1061_ sky130_fd_sc_hd__a21o_1
X_2262_ _0943_ _0948_ _0926_ VGND VGND VDPWR VDPWR _0051_ sky130_fd_sc_hd__a21oi_1
X_2193_ _0877_ _0882_ _0858_ VGND VGND VDPWR VDPWR _0048_ sky130_fd_sc_hd__a21oi_1
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[42\].clock_gate clknet_leaf_0_clk dig_ctrl_inst.latch_mem_inst.data_we\[42\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.gen_gclk\[42\]._gclk sky130_fd_sc_hd__dlclkp_1
X_1977_ _0666_ _0680_ _0681_ _0682_ VGND VGND VDPWR VDPWR _0683_ sky130_fd_sc_hd__or4_4
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[9\].clock_buffer dig_ctrl_inst.latch_mem_inst.gen_gclk\[9\]._gclk
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.gclk\[9\] sky130_fd_sc_hd__clkbuf_4
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[23\].clock_buffer dig_ctrl_inst.latch_mem_inst.gen_gclk\[23\]._gclk
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.gclk\[23\] sky130_fd_sc_hd__clkbuf_4
X_2529_ dig_ctrl_inst.spi_miso_o VGND VGND VDPWR VDPWR net25 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_30_137 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_167 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
Xhold58 dig_ctrl_inst.synchronizer_port_ms_i_inst.pipe\[0\] VGND VGND VDPWR VDPWR
+ net340 sky130_fd_sc_hd__dlygate4sd3_1
Xhold69 dig_ctrl_inst.spi_data_i\[7\] VGND VGND VDPWR VDPWR net351 sky130_fd_sc_hd__dlygate4sd3_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[62\].gen_latches\[7\].p_latch net189 dig_ctrl_inst.latch_mem_inst.gclk\[62\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[62\]\[7\] sky130_fd_sc_hd__dlxtp_1
Xhold47 dig_ctrl_inst.latch_mem_inst.wdata\[3\] VGND VGND VDPWR VDPWR net329 sky130_fd_sc_hd__dlygate4sd3_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[51\].gen_latches\[5\].p_latch net202 dig_ctrl_inst.latch_mem_inst.gclk\[51\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[51\]\[5\] sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[40\].gen_latches\[3\].p_latch net216 dig_ctrl_inst.latch_mem_inst.gclk\[40\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[40\]\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_44_218 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_1831_ dig_ctrl_inst.latch_mem_inst.RAM\[30\]\[4\] net72 net64 VGND VGND VDPWR VDPWR
+ _0539_ sky130_fd_sc_hd__and3_2
XFILLER_0_32_56 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
X_1900_ dig_ctrl_inst.latch_mem_inst.RAM\[33\]\[5\] _0135_ _0604_ _0605_ _0606_ VGND
+ VGND VDPWR VDPWR _0607_ sky130_fd_sc_hd__a2111o_1
X_1762_ dig_ctrl_inst.latch_mem_inst.RAM\[41\]\[3\] net119 net92 net59 VGND VGND VDPWR
+ VDPWR _0471_ sky130_fd_sc_hd__and4_1
X_1693_ dig_ctrl_inst.latch_mem_inst.RAM\[12\]\[2\] net126 net78 VGND VGND VDPWR VDPWR
+ _0403_ sky130_fd_sc_hd__and3_2
XFILLER_0_57_31 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_2314_ net368 _0973_ _0977_ VGND VGND VDPWR VDPWR _0074_ sky130_fd_sc_hd__mux2_1
X_2176_ _0252_ _0864_ _0865_ VGND VGND VDPWR VDPWR _0866_ sky130_fd_sc_hd__o21ai_1
X_2245_ net167 _0838_ _0929_ _0931_ net170 VGND VGND VDPWR VDPWR _0932_ sky130_fd_sc_hd__a221o_1
XFILLER_0_73_41 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_23_305 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput26 net26 VGND VGND VDPWR VDPWR uio_out[6] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_1_Right_1 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[55\].gen_latches\[6\].p_latch net197 dig_ctrl_inst.latch_mem_inst.gclk\[55\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[55\]\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_34_273 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_329 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_6
Xdig_ctrl_inst.latch_mem_inst.gen_words\[44\].gen_latches\[4\].p_latch net209 dig_ctrl_inst.latch_mem_inst.gclk\[44\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[44\]\[4\] sky130_fd_sc_hd__dlxtp_1
X_2030_ dig_ctrl_inst.latch_mem_inst.RAM\[43\]\[7\] _0143_ _0696_ _0697_ _0707_ VGND
+ VGND VDPWR VDPWR _0735_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_43_77 VDPWR VGND VDPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_55 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[33\].gen_latches\[2\].p_latch net231 dig_ctrl_inst.latch_mem_inst.gclk\[33\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[33\]\[2\] sky130_fd_sc_hd__dlxtp_1
X_1745_ dig_ctrl_inst.latch_mem_inst.RAM\[63\]\[3\] _0160_ _0277_ dig_ctrl_inst.latch_mem_inst.RAM\[4\]\[3\]
+ VGND VGND VDPWR VDPWR _0454_ sky130_fd_sc_hd__a22o_1
X_1814_ dig_ctrl_inst.latch_mem_inst.RAM\[60\]\[4\] net76 net45 VGND VGND VDPWR VDPWR
+ _0522_ sky130_fd_sc_hd__and3_2
XFILLER_0_68_85 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_8
Xdig_ctrl_inst.latch_mem_inst.gen_words\[22\].gen_latches\[0\].p_latch net245 dig_ctrl_inst.latch_mem_inst.gclk\[22\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[22\]\[0\] sky130_fd_sc_hd__dlxtp_1
X_1676_ dig_ctrl_inst.latch_mem_inst.RAM\[35\]\[1\] _0137_ _0353_ _0356_ _0368_ VGND
+ VGND VDPWR VDPWR _0387_ sky130_fd_sc_hd__a2111o_1
X_2159_ _0247_ _0849_ _0787_ _0248_ VGND VGND VDPWR VDPWR _0850_ sky130_fd_sc_hd__o2bb2a_1
X_2228_ net138 _0783_ _0915_ VGND VGND VDPWR VDPWR _0916_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_63_335 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_39_Left_117 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_287 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[59\].gen_latches\[7\].p_latch net188 dig_ctrl_inst.latch_mem_inst.gclk\[59\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[59\]\[7\] sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[10\].gen_latches\[7\].p_latch net185 dig_ctrl_inst.latch_mem_inst.gclk\[10\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[10\]\[7\] sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_48_Left_126 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[4\].gen_latches\[0\].p_latch net246 dig_ctrl_inst.latch_mem_inst.gclk\[4\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[4\]\[0\] sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_57_Left_135 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[48\].gen_latches\[5\].p_latch net201 dig_ctrl_inst.latch_mem_inst.gclk\[48\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[48\]\[5\] sky130_fd_sc_hd__dlxtp_1
X_1461_ _1003_ _1096_ _0189_ _0184_ VGND VGND VDPWR VDPWR _0192_ sky130_fd_sc_hd__o31a_1
X_1530_ _1103_ net160 VGND VGND VDPWR VDPWR _0243_ sky130_fd_sc_hd__nor2_1
X_1392_ net149 _0151_ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.data_we\[53\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_22_287 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_2013_ dig_ctrl_inst.latch_mem_inst.RAM\[19\]\[7\] _0122_ _0156_ dig_ctrl_inst.latch_mem_inst.RAM\[59\]\[7\]
+ VGND VGND VDPWR VDPWR _0718_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_66_Left_144 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[37\].gen_latches\[3\].p_latch net217 dig_ctrl_inst.latch_mem_inst.gclk\[37\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[37\]\[3\] sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_75_Left_153 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_15_clk clknet_1_0__leaf_clk VGND VGND VDPWR VDPWR clknet_leaf_15_clk
+ sky130_fd_sc_hd__clkbuf_8
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[16\].clock_buffer dig_ctrl_inst.latch_mem_inst.gen_gclk\[16\]._gclk
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.gclk\[16\] sky130_fd_sc_hd__clkbuf_4
Xhold100 dig_ctrl_inst.spi_addr\[0\] VGND VGND VDPWR VDPWR net382 sky130_fd_sc_hd__dlygate4sd3_1
X_1728_ dig_ctrl_inst.latch_mem_inst.RAM\[41\]\[2\] _0141_ _0406_ _0408_ _0412_ VGND
+ VGND VDPWR VDPWR _0438_ sky130_fd_sc_hd__a2111o_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[26\].gen_latches\[1\].p_latch net236 dig_ctrl_inst.latch_mem_inst.gclk\[26\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[26\]\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_0_181 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_6
X_1659_ dig_ctrl_inst.latch_mem_inst.RAM\[44\]\[1\] net76 net54 VGND VGND VDPWR VDPWR
+ _0370_ sky130_fd_sc_hd__and3_2
XTAP_TAPCELL_ROW_56_503 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2524__273 VGND VGND VDPWR VDPWR _2524__273/HI net273 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_4_191 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2531__277 VGND VGND VDPWR VDPWR _2531__277/HI net277 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_62_539 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_151 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[8\].gen_latches\[1\].p_latch net235 dig_ctrl_inst.latch_mem_inst.gclk\[8\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[8\]\[1\] sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_70_583 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_34 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_6
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[47\].clock_gate clknet_leaf_18_clk dig_ctrl_inst.latch_mem_inst.data_we\[47\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.gen_gclk\[47\]._gclk sky130_fd_sc_hd__dlclkp_1
X_1444_ dig_ctrl_inst.spi_receiver_inst.spi_cs_sync dig_ctrl_inst.spi_receiver_inst.spi_sclk_sync
+ dig_ctrl_inst.spi_receiver_inst.spi_sclk_delayed VGND VGND VDPWR VDPWR _0180_ sky130_fd_sc_hd__or3b_4
Xclkbuf_leaf_4_clk clknet_1_1__leaf_clk VGND VGND VDPWR VDPWR clknet_leaf_4_clk sky130_fd_sc_hd__clkbuf_8
X_2493_ clknet_leaf_6_clk _0092_ net179 VGND VGND VDPWR VDPWR dig_ctrl_inst.spi_data_i\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_1375_ net78 net58 VGND VGND VDPWR VDPWR _0144_ sky130_fd_sc_hd__and2_1
X_1513_ _0998_ dig_ctrl_inst.cpu_inst.r2\[6\] dig_ctrl_inst.cpu_inst.r1\[6\] _1022_
+ net299 VGND VGND VDPWR VDPWR _0226_ sky130_fd_sc_hd__a221o_1
XFILLER_0_10_279 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_8
X_1159__1 clknet_leaf_4_clk VGND VGND VDPWR VDPWR net282 sky130_fd_sc_hd__inv_2
XFILLER_0_45_165 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_327 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_240 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_271 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_313 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[19\].gen_latches\[0\].p_latch net244 dig_ctrl_inst.latch_mem_inst.gclk\[19\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[19\]\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_5_262 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_1_172 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout83 net84 VGND VGND VDPWR VDPWR net83 sky130_fd_sc_hd__buf_2
Xfanout50 _0147_ VGND VGND VDPWR VDPWR net50 sky130_fd_sc_hd__buf_4
Xfanout94 net95 VGND VGND VDPWR VDPWR net94 sky130_fd_sc_hd__buf_1
XFILLER_0_10_48 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
Xfanout61 net67 VGND VGND VDPWR VDPWR net61 sky130_fd_sc_hd__clkbuf_2
Xfanout72 net75 VGND VGND VDPWR VDPWR net72 sky130_fd_sc_hd__clkbuf_4
X_1160_ _1002_ dig_ctrl_inst.spi_addr\[3\] VGND VGND VDPWR VDPWR _1008_ sky130_fd_sc_hd__or2_1
X_1993_ dig_ctrl_inst.latch_mem_inst.RAM\[56\]\[7\] net88 net48 VGND VGND VDPWR VDPWR
+ _0698_ sky130_fd_sc_hd__and3_2
XTAP_TAPCELL_ROW_15_252 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_209 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_85 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
X_2476_ clknet_leaf_2_clk _0082_ net172 VGND VGND VDPWR VDPWR dig_ctrl_inst.spi_data_o\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_1358_ net148 net109 net51 VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.data_we\[34\]
+ sky130_fd_sc_hd__and3_2
X_1427_ net258 net255 dig_ctrl_inst.cpu_inst.r3\[7\] VGND VGND VDPWR VDPWR _0168_
+ sky130_fd_sc_hd__and3_2
X_1289_ net304 _1078_ _1093_ VGND VGND VDPWR VDPWR _1134_ sky130_fd_sc_hd__and3_4
Xclkload3 clknet_leaf_12_clk VGND VGND VDPWR VDPWR clkload3/Y sky130_fd_sc_hd__clkinv_8
XTAP_TAPCELL_ROW_21_288 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout240 net241 VGND VGND VDPWR VDPWR net240 sky130_fd_sc_hd__clkbuf_2
Xfanout251 dig_ctrl_inst.mode_sync VGND VGND VDPWR VDPWR net251 sky130_fd_sc_hd__clkbuf_2
Xfanout262 net264 VGND VGND VDPWR VDPWR net262 sky130_fd_sc_hd__buf_4
XFILLER_0_56_238 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_205 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[62\].clock_buffer dig_ctrl_inst.latch_mem_inst.gen_gclk\[62\]._gclk
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.gclk\[62\] sky130_fd_sc_hd__clkbuf_4
X_2330_ dig_ctrl_inst.spi_data_o\[2\] dig_ctrl_inst.spi_data_o\[3\] _0180_ VGND VGND
+ VDPWR VDPWR _0082_ sky130_fd_sc_hd__mux2_1
X_2192_ _0754_ _0880_ _0881_ _0756_ net41 VGND VGND VDPWR VDPWR _0882_ sky130_fd_sc_hd__o221a_1
X_1212_ net300 _1056_ _1057_ _1058_ _1059_ VGND VGND VDPWR VDPWR _1060_ sky130_fd_sc_hd__o41a_2
XFILLER_0_46_11 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
X_2261_ _0754_ _0946_ _0947_ _0756_ net41 VGND VGND VDPWR VDPWR _0948_ sky130_fd_sc_hd__o221a_1
XFILLER_0_47_205 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[63\].gen_latches\[2\].p_latch net226 dig_ctrl_inst.latch_mem_inst.gclk\[63\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[63\]\[2\] sky130_fd_sc_hd__dlxtp_1
X_1976_ dig_ctrl_inst.latch_mem_inst.RAM\[41\]\[6\] _0141_ _0626_ _0627_ _0629_ VGND
+ VGND VDPWR VDPWR _0682_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_15_146 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
X_2528_ net275 VGND VGND VDPWR VDPWR uio_out[1] sky130_fd_sc_hd__buf_2
XFILLER_0_60_3 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_341 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
Xhold59 dig_ctrl_inst.synchronizer_port_i_inst\[0\].pipe\[0\] VGND VGND VDPWR VDPWR
+ net341 sky130_fd_sc_hd__dlygate4sd3_1
Xhold48 dig_ctrl_inst.synchronizer_port_i_inst\[3\].pipe\[0\] VGND VGND VDPWR VDPWR
+ net330 sky130_fd_sc_hd__dlygate4sd3_1
X_2459_ clknet_leaf_11_clk _0067_ net142 VGND VGND VDPWR VDPWR dig_ctrl_inst.cpu_inst.r2\[6\]
+ sky130_fd_sc_hd__dfrtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[52\].gen_latches\[0\].p_latch net241 dig_ctrl_inst.latch_mem_inst.gclk\[52\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[52\]\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_46_282 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[40\].gen_latches\[7\].p_latch net185 dig_ctrl_inst.latch_mem_inst.gclk\[40\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[40\]\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_16_69 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
X_1761_ dig_ctrl_inst.latch_mem_inst.RAM\[7\]\[3\] net126 net106 net101 VGND VGND
+ VDPWR VDPWR _0470_ sky130_fd_sc_hd__and4_1
X_1830_ _0154_ dig_ctrl_inst.latch_mem_inst.RAM\[57\]\[4\] _0535_ _0536_ _0537_ VGND
+ VGND VDPWR VDPWR _0538_ sky130_fd_sc_hd__a2111o_1
X_1692_ dig_ctrl_inst.latch_mem_inst.RAM\[56\]\[2\] net88 net50 VGND VGND VDPWR VDPWR
+ _0402_ sky130_fd_sc_hd__and3_2
X_2313_ net376 _0972_ _0977_ VGND VGND VDPWR VDPWR _0073_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_48_450 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2175_ _0252_ _0864_ _0788_ VGND VGND VDPWR VDPWR _0865_ sky130_fd_sc_hd__a21oi_1
X_2244_ _0840_ _0886_ _0930_ VGND VGND VDPWR VDPWR _0931_ sky130_fd_sc_hd__and3_2
XPHY_EDGE_ROW_11_Left_89 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
X_1959_ dig_ctrl_inst.latch_mem_inst.RAM\[37\]\[6\] _0138_ _0624_ _0647_ _0659_ VGND
+ VGND VDPWR VDPWR _0665_ sky130_fd_sc_hd__a2111o_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[56\].gen_latches\[1\].p_latch net238 dig_ctrl_inst.latch_mem_inst.gclk\[56\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[56\]\[1\] sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_31_350 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput27 net27 VGND VGND VDPWR VDPWR uio_out[7] sky130_fd_sc_hd__buf_2
Xoutput16 net16 VGND VGND VDPWR VDPWR clk_o sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_54_486 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[0\].gen_latches\[3\].p_latch net218 dig_ctrl_inst.latch_mem_inst.gclk\[0\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[0\]\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_43_89 VDPWR VGND VDPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_0_clk clk VGND VGND VDPWR VDPWR clknet_0_clk sky130_fd_sc_hd__clkbuf_16
Xdig_ctrl_inst.latch_mem_inst.gen_words\[33\].gen_latches\[6\].p_latch net192 dig_ctrl_inst.latch_mem_inst.gclk\[33\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[33\]\[6\] sky130_fd_sc_hd__dlxtp_1
X_1744_ dig_ctrl_inst.latch_mem_inst.RAM\[14\]\[3\] _0116_ _0279_ dig_ctrl_inst.latch_mem_inst.RAM\[6\]\[3\]
+ _0452_ VGND VGND VDPWR VDPWR _0453_ sky130_fd_sc_hd__a221o_1
XFILLER_0_4_179 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
X_1813_ dig_ctrl_inst.latch_mem_inst.RAM\[44\]\[4\] net76 net54 VGND VGND VDPWR VDPWR
+ _0521_ sky130_fd_sc_hd__and3_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[22\].gen_latches\[4\].p_latch net212 dig_ctrl_inst.latch_mem_inst.gclk\[22\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[22\]\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_0_341 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_1675_ _0379_ _0380_ _0381_ _0385_ VGND VGND VDPWR VDPWR _0386_ sky130_fd_sc_hd__or4_1
XPHY_EDGE_ROW_15_Right_15 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
X_2158_ net167 _0790_ _0785_ VGND VGND VDPWR VDPWR _0849_ sky130_fd_sc_hd__a21bo_1
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[54\].clock_gate clknet_leaf_16_clk dig_ctrl_inst.latch_mem_inst.data_we\[54\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.gen_gclk\[54\]._gclk sky130_fd_sc_hd__dlclkp_1
X_2089_ net168 _0781_ _0774_ net171 VGND VGND VDPWR VDPWR _0782_ sky130_fd_sc_hd__a211o_1
X_2227_ dig_ctrl_inst.cpu_inst.data\[5\] _0743_ _0825_ net159 VGND VGND VDPWR VDPWR
+ _0915_ sky130_fd_sc_hd__a22o_1
XFILLER_0_23_3 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_24_Right_24 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[11\].gen_latches\[2\].p_latch net229 dig_ctrl_inst.latch_mem_inst.gclk\[11\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[11\]\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_48_333 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_33_Right_33 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[49\].gen_latches\[0\].p_latch net244 dig_ctrl_inst.latch_mem_inst.gclk\[49\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[49\]\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_66_141 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_42_Right_42 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_51_Right_51 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[4\].gen_latches\[4\].p_latch net213 dig_ctrl_inst.latch_mem_inst.gclk\[4\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[4\]\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_1_105 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[55\].clock_buffer dig_ctrl_inst.latch_mem_inst.gen_gclk\[55\]._gclk
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.gclk\[55\] sky130_fd_sc_hd__clkbuf_4
X_1460_ _1003_ _0189_ VGND VGND VDPWR VDPWR _0191_ sky130_fd_sc_hd__nor2_1
X_1391_ net117 net100 net45 VGND VGND VDPWR VDPWR _0151_ sky130_fd_sc_hd__and3_2
X_2012_ _0714_ _0715_ _0716_ VGND VGND VDPWR VDPWR _0717_ sky130_fd_sc_hd__or3_1
XPHY_EDGE_ROW_60_Right_60 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_44 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[37\].gen_latches\[7\].p_latch net186 dig_ctrl_inst.latch_mem_inst.gclk\[37\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[37\]\[7\] sky130_fd_sc_hd__dlxtp_1
Xhold101 net23 VGND VGND VDPWR VDPWR net383 sky130_fd_sc_hd__dlygate4sd3_1
X_1727_ dig_ctrl_inst.latch_mem_inst.RAM\[39\]\[2\] _0139_ _0403_ _0407_ _0409_ VGND
+ VGND VDPWR VDPWR _0437_ sky130_fd_sc_hd__a2111o_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[26\].gen_latches\[5\].p_latch net203 dig_ctrl_inst.latch_mem_inst.gclk\[26\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[26\]\[5\] sky130_fd_sc_hd__dlxtp_1
X_1658_ dig_ctrl_inst.latch_mem_inst.RAM\[32\]\[1\] net128 net55 VGND VGND VDPWR VDPWR
+ _0369_ sky130_fd_sc_hd__and3_2
X_1589_ dig_ctrl_inst.latch_mem_inst.RAM\[14\]\[0\] net123 net74 VGND VGND VDPWR VDPWR
+ _0301_ sky130_fd_sc_hd__and3_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[15\].gen_latches\[3\].p_latch net222 dig_ctrl_inst.latch_mem_inst.gclk\[15\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[15\]\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_48_141 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_14_Left_92 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_70_584 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[8\].gen_latches\[5\].p_latch net204 dig_ctrl_inst.latch_mem_inst.gclk\[8\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[8\]\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_40_24 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
X_2492_ clknet_leaf_4_clk _0091_ net179 VGND VGND VDPWR VDPWR dig_ctrl_inst.spi_data_i\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_57 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
X_1512_ net265 net262 dig_ctrl_inst.cpu_inst.r3\[6\] VGND VGND VDPWR VDPWR _0225_
+ sky130_fd_sc_hd__and3_2
XFILLER_0_10_203 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
X_1443_ _0177_ _0178_ _0179_ _1039_ _1027_ VGND VGND VDPWR VDPWR dig_ctrl_inst.cpu_inst.stb_o
+ sky130_fd_sc_hd__o32a_1
X_1374_ net152 _0143_ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.data_we\[43\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_65_87 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_18_272 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_144 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_111 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_317 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[19\].gen_latches\[4\].p_latch net208 dig_ctrl_inst.latch_mem_inst.gclk\[19\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[19\]\[4\] sky130_fd_sc_hd__dlxtp_1
Xfanout73 net74 VGND VGND VDPWR VDPWR net73 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_1_173 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout62 net63 VGND VGND VDPWR VDPWR net62 sky130_fd_sc_hd__clkbuf_2
Xfanout51 net53 VGND VGND VDPWR VDPWR net51 sky130_fd_sc_hd__buf_4
XFILLER_0_51_125 VDPWR VGND VDPWR VGND sky130_ef_sc_hd__decap_12
Xfanout95 _1138_ VGND VGND VDPWR VDPWR net95 sky130_fd_sc_hd__buf_4
Xfanout84 _1144_ VGND VGND VDPWR VDPWR net84 sky130_fd_sc_hd__buf_4
XFILLER_0_10_27 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_339 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_57 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
Xclkload10 clknet_leaf_3_clk VGND VGND VDPWR VDPWR clkload10/Y sky130_fd_sc_hd__clkinv_4
XFILLER_0_51_34 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
X_1992_ dig_ctrl_inst.latch_mem_inst.RAM\[18\]\[7\] net111 net64 VGND VGND VDPWR VDPWR
+ _0697_ sky130_fd_sc_hd__and3_2
XTAP_TAPCELL_ROW_15_253 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2475_ clknet_leaf_4_clk _0081_ net172 VGND VGND VDPWR VDPWR dig_ctrl_inst.spi_data_o\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_1426_ net250 dig_ctrl_inst.spi_data_o\[6\] _0162_ _0167_ VGND VGND VDPWR VDPWR dig_ctrl_inst.data_out\[6\]
+ sky130_fd_sc_hd__a22o_1
X_1357_ net111 net58 VGND VGND VDPWR VDPWR _0136_ sky130_fd_sc_hd__and2_1
X_1288_ net150 net120 net109 VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.data_we\[2\]
+ sky130_fd_sc_hd__and3_2
XFILLER_0_58_291 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_21_289 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload4 clknet_leaf_13_clk VGND VGND VDPWR VDPWR clkload4/Y sky130_fd_sc_hd__clkinv_4
Xfanout230 net231 VGND VGND VDPWR VDPWR net230 sky130_fd_sc_hd__clkbuf_2
Xfanout263 net264 VGND VGND VDPWR VDPWR net263 sky130_fd_sc_hd__buf_6
Xfanout241 net242 VGND VGND VDPWR VDPWR net241 sky130_fd_sc_hd__clkbuf_2
Xfanout252 dig_ctrl_inst.cpu_inst.instr\[5\] VGND VGND VDPWR VDPWR net252 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_64_250 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[48\].clock_buffer dig_ctrl_inst.latch_mem_inst.gen_gclk\[48\]._gclk
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.gclk\[48\] sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_12_234 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_15 VDPWR VGND VDPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_191 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_309 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_6
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[59\].clock_gate clknet_leaf_0_clk dig_ctrl_inst.latch_mem_inst.data_we\[59\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.gen_gclk\[59\]._gclk sky130_fd_sc_hd__dlclkp_1
X_2191_ dig_ctrl_inst.synchronizer_port_i_inst\[3\].out _0802_ _0804_ dig_ctrl_inst.spi_data_o\[3\]
+ VGND VGND VDPWR VDPWR _0881_ sky130_fd_sc_hd__a22oi_1
X_2260_ dig_ctrl_inst.synchronizer_port_i_inst\[6\].out _0802_ _0804_ dig_ctrl_inst.spi_data_o\[6\]
+ VGND VGND VDPWR VDPWR _0947_ sky130_fd_sc_hd__a22oi_2
X_1211_ net268 net263 dig_ctrl_inst.cpu_inst.r0\[2\] VGND VGND VDPWR VDPWR _1059_
+ sky130_fd_sc_hd__or3_1
XFILLER_0_46_67 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_66 VDPWR VGND VDPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_242 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[63\].gen_latches\[6\].p_latch net194 dig_ctrl_inst.latch_mem_inst.gclk\[63\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[63\]\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_11_81 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_169 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
X_1975_ dig_ctrl_inst.latch_mem_inst.RAM\[51\]\[6\] _0149_ _0628_ _0631_ _0653_ VGND
+ VGND VDPWR VDPWR _0681_ sky130_fd_sc_hd__a2111o_1
X_1409_ net153 net73 net48 VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.data_we\[62\]
+ sky130_fd_sc_hd__and3_2
X_2527_ net274 VGND VGND VDPWR VDPWR uio_out[0] sky130_fd_sc_hd__buf_2
X_2458_ clknet_leaf_7_clk _0066_ net143 VGND VGND VDPWR VDPWR dig_ctrl_inst.cpu_inst.r2\[5\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold49 dig_ctrl_inst.synchronizer_port_i_inst\[5\].pipe\[0\] VGND VGND VDPWR VDPWR
+ net331 sky130_fd_sc_hd__dlygate4sd3_1
X_2389_ clknet_leaf_4_clk net334 net172 VGND VGND VDPWR VDPWR dig_ctrl_inst.synchronizer_port_i_inst\[2\].out
+ sky130_fd_sc_hd__dfrtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[52\].gen_latches\[4\].p_latch net209 dig_ctrl_inst.latch_mem_inst.gclk\[52\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[52\]\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_46_250 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_34_370 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[61\].clock_gate clknet_leaf_15_clk dig_ctrl_inst.latch_mem_inst.data_we\[61\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.gen_gclk\[61\]._gclk sky130_fd_sc_hd__dlclkp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[41\].gen_latches\[2\].p_latch net225 dig_ctrl_inst.latch_mem_inst.gclk\[41\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[41\]\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_21_106 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_6
Xdig_ctrl_inst.latch_mem_inst.gen_words\[30\].gen_latches\[0\].p_latch net244 dig_ctrl_inst.latch_mem_inst.gclk\[30\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[30\]\[0\] sky130_fd_sc_hd__dlxtp_1
X_1691_ dig_ctrl_inst.latch_mem_inst.RAM\[15\]\[2\] net127 net106 net82 VGND VGND
+ VDPWR VDPWR _0401_ sky130_fd_sc_hd__and4_1
XFILLER_0_52_253 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_242 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_328 VDPWR VGND VDPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_2_Left_80 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
X_1760_ _0466_ _0467_ _0468_ VGND VGND VDPWR VDPWR _0469_ sky130_fd_sc_hd__or3_1
X_2312_ net370 _0971_ _0977_ VGND VGND VDPWR VDPWR _0072_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_48_451 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2174_ _0248_ _0852_ _0246_ VGND VGND VDPWR VDPWR _0864_ sky130_fd_sc_hd__o21a_1
X_2243_ net158 _0775_ _0778_ _0770_ VGND VGND VDPWR VDPWR _0930_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_31_351 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_250 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_133 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
Xoutput17 net17 VGND VGND VDPWR VDPWR port_ms_o[0] sky130_fd_sc_hd__buf_2
Xoutput28 net28 VGND VGND VDPWR VDPWR uo_out[0] sky130_fd_sc_hd__buf_2
X_1958_ _0640_ _0652_ _0654_ _0655_ VGND VGND VDPWR VDPWR _0664_ sky130_fd_sc_hd__or4_1
X_1889_ dig_ctrl_inst.latch_mem_inst.RAM\[43\]\[5\] _0143_ _0149_ dig_ctrl_inst.latch_mem_inst.RAM\[51\]\[5\]
+ VGND VGND VDPWR VDPWR _0596_ sky130_fd_sc_hd__a22o_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[56\].gen_latches\[5\].p_latch net204 dig_ctrl_inst.latch_mem_inst.gclk\[56\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[56\]\[5\] sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[5\].clock_buffer dig_ctrl_inst.latch_mem_inst.gen_gclk\[5\]._gclk
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.gclk\[5\] sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_54_487 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[45\].gen_latches\[3\].p_latch net219 dig_ctrl_inst.latch_mem_inst.gclk\[45\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[45\]\[3\] sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[34\].gen_latches\[1\].p_latch net233 dig_ctrl_inst.latch_mem_inst.gclk\[34\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[34\]\[1\] sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[0\].gen_latches\[7\].p_latch net190 dig_ctrl_inst.latch_mem_inst.gclk\[0\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[0\]\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_27_69 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_45_432 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1743_ dig_ctrl_inst.latch_mem_inst.RAM\[1\]\[3\] _1130_ _0123_ dig_ctrl_inst.latch_mem_inst.RAM\[20\]\[3\]
+ VGND VGND VDPWR VDPWR _0452_ sky130_fd_sc_hd__a22o_1
X_1674_ dig_ctrl_inst.latch_mem_inst.RAM\[57\]\[1\] _0154_ _0355_ _0363_ _0366_ VGND
+ VGND VDPWR VDPWR _0385_ sky130_fd_sc_hd__a2111o_1
X_1812_ dig_ctrl_inst.latch_mem_inst.RAM\[16\]\[4\] net129 net64 VGND VGND VDPWR VDPWR
+ _0520_ sky130_fd_sc_hd__and3_2
X_2226_ _0243_ _0785_ _0793_ _0242_ _0913_ VGND VGND VDPWR VDPWR _0914_ sky130_fd_sc_hd__o221a_1
X_2157_ _0246_ _0793_ _0847_ VGND VGND VDPWR VDPWR _0848_ sky130_fd_sc_hd__o21ba_1
X_2088_ _0768_ _0777_ _0780_ _0765_ VGND VGND VDPWR VDPWR _0781_ sky130_fd_sc_hd__o22a_1
XFILLER_0_16_3 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_153 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_337 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_51_468 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_231 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_253 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[11\].gen_latches\[6\].p_latch net195 dig_ctrl_inst.latch_mem_inst.gclk\[11\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[11\]\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_31_278 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[49\].gen_latches\[4\].p_latch net212 dig_ctrl_inst.latch_mem_inst.gclk\[49\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[49\]\[4\] sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[38\].gen_latches\[2\].p_latch net228 dig_ctrl_inst.latch_mem_inst.gclk\[38\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[38\]\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_1_139 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
X_1390_ net151 net96 net43 VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.data_we\[52\]
+ sky130_fd_sc_hd__and3_2
X_2011_ dig_ctrl_inst.latch_mem_inst.RAM\[7\]\[7\] _1139_ _0117_ dig_ctrl_inst.latch_mem_inst.RAM\[15\]\[7\]
+ VGND VGND VDPWR VDPWR _0716_ sky130_fd_sc_hd__a22o_1
XFILLER_0_49_109 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[27\].gen_latches\[0\].p_latch net241 dig_ctrl_inst.latch_mem_inst.gclk\[27\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[27\]\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_70_99 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XFILLER_0_70_11 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_307 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_1726_ dig_ctrl_inst.latch_mem_inst.RAM\[11\]\[2\] _1145_ _0399_ _0401_ _0410_ VGND
+ VGND VDPWR VDPWR _0436_ sky130_fd_sc_hd__a2111o_1
X_1657_ dig_ctrl_inst.latch_mem_inst.RAM\[8\]\[1\] net121 net86 VGND VGND VDPWR VDPWR
+ _0368_ sky130_fd_sc_hd__and3_2
XFILLER_0_13_289 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
Xhold102 dig_ctrl_inst.cpu_inst.r2\[7\] VGND VGND VDPWR VDPWR net384 sky130_fd_sc_hd__dlygate4sd3_1
X_1588_ dig_ctrl_inst.latch_mem_inst.RAM\[48\]\[0\] net130 net45 VGND VGND VDPWR VDPWR
+ _0300_ sky130_fd_sc_hd__and3_2
XFILLER_0_0_194 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
X_2209_ _0239_ _0785_ _0895_ _0897_ VGND VGND VDPWR VDPWR _0898_ sky130_fd_sc_hd__o211a_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[15\].gen_latches\[7\].p_latch net189 dig_ctrl_inst.latch_mem_inst.gclk\[15\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[15\]\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_48_175 VDPWR VGND VDPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_167 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_197 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_272 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[9\].gen_latches\[0\].p_latch net241 dig_ctrl_inst.latch_mem_inst.gclk\[9\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[9\]\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_5_3 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_70_585 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_337 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
X_2491_ clknet_leaf_5_clk _0090_ net178 VGND VGND VDPWR VDPWR dig_ctrl_inst.spi_data_i\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_1442_ dig_ctrl_inst.cpu_inst.cpu_state\[1\] dig_ctrl_inst.cpu_inst.prev_state\[1\]
+ VGND VGND VDPWR VDPWR _0179_ sky130_fd_sc_hd__xor2_1
X_1511_ _1006_ _0220_ _0224_ _0204_ VGND VGND VDPWR VDPWR _0024_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_65_55 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_1373_ net108 net92 net59 VGND VGND VDPWR VDPWR _0143_ sky130_fd_sc_hd__and3_2
XTAP_TAPCELL_ROW_61_530 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_81 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_18_273 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_231 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[12\].clock_buffer dig_ctrl_inst.latch_mem_inst.gen_gclk\[12\]._gclk
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.gclk\[12\] sky130_fd_sc_hd__clkbuf_4
X_1709_ dig_ctrl_inst.latch_mem_inst.RAM\[1\]\[2\] _1130_ _0160_ dig_ctrl_inst.latch_mem_inst.RAM\[63\]\[2\]
+ _0418_ VGND VGND VDPWR VDPWR _0419_ sky130_fd_sc_hd__a221o_1
Xfanout74 net75 VGND VGND VDPWR VDPWR net74 sky130_fd_sc_hd__buf_4
Xfanout41 _0758_ VGND VGND VDPWR VDPWR net41 sky130_fd_sc_hd__buf_2
XFILLER_0_36_167 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
Xfanout96 net98 VGND VGND VDPWR VDPWR net96 sky130_fd_sc_hd__buf_2
Xfanout52 net53 VGND VGND VDPWR VDPWR net52 sky130_fd_sc_hd__clkbuf_2
Xfanout63 net67 VGND VGND VDPWR VDPWR net63 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_51_137 VDPWR VGND VDPWR VGND sky130_ef_sc_hd__decap_12
Xdig_ctrl_inst.latch_mem_inst.gen_words\[60\].gen_latches\[0\].p_latch net244 dig_ctrl_inst.latch_mem_inst.gclk\[60\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[60\]\[0\] sky130_fd_sc_hd__dlxtp_1
Xclkload11 clknet_leaf_4_clk VGND VGND VDPWR VDPWR clkload11/Y sky130_fd_sc_hd__bufinv_16
XTAP_TAPCELL_ROW_15_254 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1991_ dig_ctrl_inst.latch_mem_inst.RAM\[16\]\[7\] net130 net64 VGND VGND VDPWR VDPWR
+ _0696_ sky130_fd_sc_hd__and3_2
XFILLER_0_76_43 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
X_2474_ clknet_leaf_4_clk _0080_ net172 VGND VGND VDPWR VDPWR dig_ctrl_inst.spi_data_o\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_1425_ _1018_ _0163_ _0164_ _0165_ _0166_ VGND VGND VDPWR VDPWR _0167_ sky130_fd_sc_hd__o41a_4
XFILLER_0_2_278 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_1287_ net120 net110 VGND VGND VDPWR VDPWR _1133_ sky130_fd_sc_hd__and2_2
X_1356_ net150 _0135_ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.data_we\[33\]
+ sky130_fd_sc_hd__and2_1
Xclkload5 clknet_leaf_15_clk VGND VGND VDPWR VDPWR clkload5/Y sky130_fd_sc_hd__inv_8
Xfanout231 net324 VGND VGND VDPWR VDPWR net231 sky130_fd_sc_hd__buf_2
Xfanout220 net221 VGND VGND VDPWR VDPWR net220 sky130_fd_sc_hd__clkbuf_2
Xfanout264 dig_ctrl_inst.cpu_inst.arg0\[1\] VGND VGND VDPWR VDPWR net264 sky130_fd_sc_hd__buf_4
Xfanout242 net247 VGND VGND VDPWR VDPWR net242 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_6_200 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout253 dig_ctrl_inst.cpu_inst.instr\[4\] VGND VGND VDPWR VDPWR net253 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_12_235 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_27 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_12 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
X_2190_ _0878_ _0879_ VGND VGND VDPWR VDPWR _0880_ sky130_fd_sc_hd__nand2b_1
X_1210_ net263 dig_ctrl_inst.cpu_inst.r1\[2\] VGND VGND VDPWR VDPWR _1058_ sky130_fd_sc_hd__and2b_1
XFILLER_0_1_15 VDPWR VGND VDPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_78 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_6
X_1974_ dig_ctrl_inst.latch_mem_inst.RAM\[53\]\[6\] _0151_ _0634_ _0645_ _0651_ VGND
+ VGND VDPWR VDPWR _0680_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_7_337 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
X_2526_ net281 VGND VGND VDPWR VDPWR uio_oe[7] sky130_fd_sc_hd__buf_2
X_1408_ net73 net49 VGND VGND VDPWR VDPWR _0159_ sky130_fd_sc_hd__and2_2
X_2388_ clknet_leaf_4_clk net5 net174 VGND VGND VDPWR VDPWR dig_ctrl_inst.synchronizer_port_i_inst\[2\].pipe\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_46_3 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_8
X_2457_ clknet_leaf_7_clk _0065_ net143 VGND VGND VDPWR VDPWR dig_ctrl_inst.cpu_inst.r2\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_1339_ net149 net86 net67 VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.data_we\[24\]
+ sky130_fd_sc_hd__and3_2
XTAP_TAPCELL_ROW_34_371 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[41\].gen_latches\[6\].p_latch net193 dig_ctrl_inst.latch_mem_inst.gclk\[41\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[41\]\[6\] sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[30\].gen_latches\[4\].p_latch net209 dig_ctrl_inst.latch_mem_inst.gclk\[30\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[30\]\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_32_15 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
X_1690_ dig_ctrl_inst.latch_mem_inst.RAM\[38\]\[2\] net95 net58 VGND VGND VDPWR VDPWR
+ _0400_ sky130_fd_sc_hd__and3_2
X_2311_ net373 _0970_ _0977_ VGND VGND VDPWR VDPWR _0071_ sky130_fd_sc_hd__mux2_1
X_2242_ _0836_ _0887_ VGND VGND VDPWR VDPWR _0929_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_48_452 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2173_ _0772_ _0860_ _0861_ _0862_ net170 VGND VGND VDPWR VDPWR _0863_ sky130_fd_sc_hd__a311o_1
X_1957_ dig_ctrl_inst.latch_mem_inst.RAM\[7\]\[6\] _1139_ _0157_ dig_ctrl_inst.latch_mem_inst.RAM\[60\]\[6\]
+ VGND VGND VDPWR VDPWR _0663_ sky130_fd_sc_hd__a22o_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[57\].gen_latches\[0\].p_latch net245 dig_ctrl_inst.latch_mem_inst.gclk\[57\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[57\]\[0\] sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_31_352 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_262 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
Xoutput29 net29 VGND VGND VDPWR VDPWR uo_out[1] sky130_fd_sc_hd__buf_2
X_2509_ clknet_leaf_5_clk _0106_ net178 VGND VGND VDPWR VDPWR net20 sky130_fd_sc_hd__dfrtp_1
Xoutput18 net18 VGND VGND VDPWR VDPWR port_ms_o[1] sky130_fd_sc_hd__buf_2
X_1888_ dig_ctrl_inst.latch_mem_inst.RAM\[17\]\[5\] _0120_ _0124_ dig_ctrl_inst.latch_mem_inst.RAM\[21\]\[5\]
+ VGND VGND VDPWR VDPWR _0595_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_54_488 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[1\].gen_latches\[2\].p_latch net226 dig_ctrl_inst.latch_mem_inst.gclk\[1\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[1\]\[2\] sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[45\].gen_latches\[7\].p_latch net184 dig_ctrl_inst.latch_mem_inst.gclk\[45\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[45\]\[7\] sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_45_433 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[34\].gen_latches\[5\].p_latch net199 dig_ctrl_inst.latch_mem_inst.gclk\[34\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[34\]\[5\] sky130_fd_sc_hd__dlxtp_1
X_1811_ _0287_ _0508_ _0511_ _0518_ VGND VGND VDPWR VDPWR _0519_ sky130_fd_sc_hd__or4_1
XFILLER_0_25_210 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
XFILLER_0_68_44 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
X_1673_ _0374_ _0376_ _0382_ _0383_ VGND VGND VDPWR VDPWR _0384_ sky130_fd_sc_hd__or4_1
X_1742_ dig_ctrl_inst.latch_mem_inst.RAM\[3\]\[3\] _1135_ _0154_ dig_ctrl_inst.latch_mem_inst.RAM\[57\]\[3\]
+ _0450_ VGND VGND VDPWR VDPWR _0451_ sky130_fd_sc_hd__a221o_1
XFILLER_0_0_321 VDPWR VGND VDPWR VGND sky130_ef_sc_hd__decap_12
Xdig_ctrl_inst.latch_mem_inst.gen_words\[23\].gen_latches\[3\].p_latch net215 dig_ctrl_inst.latch_mem_inst.gclk\[23\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[23\]\[3\] sky130_fd_sc_hd__dlxtp_1
X_2225_ _0786_ _0791_ _1103_ VGND VGND VDPWR VDPWR _0913_ sky130_fd_sc_hd__mux2_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[12\].gen_latches\[1\].p_latch net237 dig_ctrl_inst.latch_mem_inst.gclk\[12\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[12\]\[1\] sky130_fd_sc_hd__dlxtp_1
Xclkbuf_leaf_18_clk clknet_1_0__leaf_clk VGND VGND VDPWR VDPWR clknet_leaf_18_clk
+ sky130_fd_sc_hd__clkbuf_8
XPHY_EDGE_ROW_5_Right_5 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
X_2087_ net157 _0779_ _0778_ VGND VGND VDPWR VDPWR _0780_ sky130_fd_sc_hd__a21o_1
X_2156_ dig_ctrl_inst.cpu_inst.data\[2\] _0743_ _0825_ net161 _0846_ VGND VGND VDPWR
+ VDPWR _0847_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_51_469 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_202 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_7 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[5\].gen_latches\[3\].p_latch net223 dig_ctrl_inst.latch_mem_inst.gclk\[5\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[5\]\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_66_176 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_338 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_42_414 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_26_Left_104 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
X_2010_ dig_ctrl_inst.latch_mem_inst.RAM\[5\]\[7\] _0278_ _0690_ _0702_ _0708_ VGND
+ VGND VDPWR VDPWR _0715_ sky130_fd_sc_hd__a2111o_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[38\].gen_latches\[6\].p_latch net195 dig_ctrl_inst.latch_mem_inst.gclk\[38\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[38\]\[6\] sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_35_Left_113 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[27\].gen_latches\[4\].p_latch net212 dig_ctrl_inst.latch_mem_inst.gclk\[27\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[27\]\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_45_327 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_44_Left_122 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
X_1725_ _0426_ _0427_ _0429_ _0431_ VGND VGND VDPWR VDPWR _0435_ sky130_fd_sc_hd__or4_1
Xhold103 net19 VGND VGND VDPWR VDPWR net385 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_7_clk clknet_1_1__leaf_clk VGND VGND VDPWR VDPWR clknet_leaf_7_clk sky130_fd_sc_hd__clkbuf_8
X_1587_ dig_ctrl_inst.latch_mem_inst.RAM\[63\]\[0\] net105 net81 net46 VGND VGND VDPWR
+ VDPWR _0299_ sky130_fd_sc_hd__and4_1
X_1656_ dig_ctrl_inst.latch_mem_inst.RAM\[30\]\[1\] net72 net64 VGND VGND VDPWR VDPWR
+ _0367_ sky130_fd_sc_hd__and3_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[16\].gen_latches\[2\].p_latch net225 dig_ctrl_inst.latch_mem_inst.gclk\[16\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[16\]\[2\] sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_53_Left_131 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_91 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_6
X_2208_ _1118_ _0786_ _0787_ _0240_ _0896_ VGND VGND VDPWR VDPWR _0897_ sky130_fd_sc_hd__o221a_1
X_2139_ _0750_ _0748_ _0830_ VGND VGND VDPWR VDPWR _0831_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_64_550 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_187 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_338 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_190 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_62_Left_140 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[9\].gen_latches\[4\].p_latch net212 dig_ctrl_inst.latch_mem_inst.gclk\[9\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[9\]\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_39_143 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_27 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_70_586 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_157 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_2490_ clknet_leaf_5_clk _0089_ net178 VGND VGND VDPWR VDPWR dig_ctrl_inst.spi_data_i\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_49_35 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_6
X_1441_ net248 _1007_ dig_ctrl_inst.cpu_inst.prev_state\[2\] _0999_ VGND VGND VDPWR
+ VDPWR _0178_ sky130_fd_sc_hd__o22ai_1
X_1510_ _1005_ _1006_ _0216_ _0223_ _0174_ VGND VGND VDPWR VDPWR _0224_ sky130_fd_sc_hd__o32a_1
X_1372_ net153 net83 net57 VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.data_we\[42\]
+ sky130_fd_sc_hd__and3_2
XFILLER_0_65_23 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_61_531 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[51\].clock_buffer dig_ctrl_inst.latch_mem_inst.gen_gclk\[51\]._gclk
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.gclk\[51\] sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_18_274 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_338 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
XFILLER_0_76_3 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_138 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_341 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_1708_ dig_ctrl_inst.latch_mem_inst.RAM\[18\]\[2\] _0121_ _0125_ dig_ctrl_inst.latch_mem_inst.RAM\[22\]\[2\]
+ VGND VGND VDPWR VDPWR _0418_ sky130_fd_sc_hd__a22o_1
XFILLER_0_30_70 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_298 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_6
X_1639_ dig_ctrl_inst.latch_mem_inst.RAM\[52\]\[1\] net96 net46 VGND VGND VDPWR VDPWR
+ _0350_ sky130_fd_sc_hd__and3_2
Xfanout97 net98 VGND VGND VDPWR VDPWR net97 sky130_fd_sc_hd__buf_2
Xfanout75 _0115_ VGND VGND VDPWR VDPWR net75 sky130_fd_sc_hd__clkbuf_2
Xfanout64 net66 VGND VGND VDPWR VDPWR net64 sky130_fd_sc_hd__buf_2
Xfanout86 net87 VGND VGND VDPWR VDPWR net86 sky130_fd_sc_hd__buf_2
Xfanout53 net54 VGND VGND VDPWR VDPWR net53 sky130_fd_sc_hd__buf_4
Xfanout42 net47 VGND VGND VDPWR VDPWR net42 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_51_149 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_9_220 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_612 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_69 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_113 VDPWR VGND VDPWR VGND sky130_ef_sc_hd__decap_12
X_1990_ dig_ctrl_inst.latch_mem_inst.RAM\[22\]\[7\] net93 net61 VGND VGND VDPWR VDPWR
+ _0695_ sky130_fd_sc_hd__and3_2
XTAP_TAPCELL_ROW_15_255 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload12 clknet_leaf_5_clk VGND VGND VDPWR VDPWR clkload12/Y sky130_fd_sc_hd__inv_8
XFILLER_0_15_319 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[60\].gen_latches\[4\].p_latch net209 dig_ctrl_inst.latch_mem_inst.gclk\[60\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[60\]\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_23_341 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_2473_ clknet_leaf_4_clk _0079_ net174 VGND VGND VDPWR VDPWR dig_ctrl_inst.spi_data_o\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_50_193 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
X_1424_ net259 net255 dig_ctrl_inst.cpu_inst.r0\[6\] VGND VGND VDPWR VDPWR _0166_
+ sky130_fd_sc_hd__or3_1
X_1355_ net131 net116 net55 VGND VGND VDPWR VDPWR _0135_ sky130_fd_sc_hd__and3_2
X_1286_ net304 _1078_ net134 net135 _1047_ VGND VGND VDPWR VDPWR _1132_ sky130_fd_sc_hd__a2111oi_1
Xclkload6 clknet_leaf_16_clk VGND VGND VDPWR VDPWR clkload6/Y sky130_fd_sc_hd__inv_6
XFILLER_0_41_193 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_6_201 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2521__279 VGND VGND VDPWR VDPWR net279 _2521__279/LO sky130_fd_sc_hd__conb_1
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[12\].clock_gate clknet_leaf_0_clk dig_ctrl_inst.latch_mem_inst.data_we\[12\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.gen_gclk\[12\]._gclk sky130_fd_sc_hd__dlclkp_1
Xfanout243 net244 VGND VGND VDPWR VDPWR net243 sky130_fd_sc_hd__clkbuf_2
Xfanout221 net223 VGND VGND VDPWR VDPWR net221 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout265 net266 VGND VGND VDPWR VDPWR net265 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_29_336 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout254 net255 VGND VGND VDPWR VDPWR net254 sky130_fd_sc_hd__buf_4
XFILLER_0_5_91 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
Xfanout210 net323 VGND VGND VDPWR VDPWR net210 sky130_fd_sc_hd__clkbuf_2
Xfanout232 net233 VGND VGND VDPWR VDPWR net232 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_12_236 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_138 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_47 VDPWR VGND VDPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_27 VDPWR VGND VDPWR VGND sky130_ef_sc_hd__decap_12
X_1973_ _0675_ _0676_ _0677_ _0678_ VGND VGND VDPWR VDPWR _0679_ sky130_fd_sc_hd__or4_4
X_2525_ net280 VGND VGND VDPWR VDPWR uio_oe[6] sky130_fd_sc_hd__buf_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[53\].gen_latches\[3\].p_latch net216 dig_ctrl_inst.latch_mem_inst.gclk\[53\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[53\]\[3\] sky130_fd_sc_hd__dlxtp_1
X_2387_ clknet_leaf_4_clk net330 net175 VGND VGND VDPWR VDPWR dig_ctrl_inst.synchronizer_port_i_inst\[3\].out
+ sky130_fd_sc_hd__dfrtp_1
X_2456_ clknet_leaf_6_clk _0064_ net145 VGND VGND VDPWR VDPWR dig_ctrl_inst.cpu_inst.r2\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_39_3 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_8
X_1338_ net86 net64 VGND VGND VDPWR VDPWR _0127_ sky130_fd_sc_hd__and2_1
X_1407_ net150 _0158_ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.data_we\[61\]
+ sky130_fd_sc_hd__and2_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[42\].gen_latches\[1\].p_latch net237 dig_ctrl_inst.latch_mem_inst.gclk\[42\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[42\]\[1\] sky130_fd_sc_hd__dlxtp_1
X_1269_ net260 net256 dig_ctrl_inst.cpu_inst.r0\[4\] VGND VGND VDPWR VDPWR _1117_
+ sky130_fd_sc_hd__or3_1
XFILLER_0_16_17 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[44\].clock_buffer dig_ctrl_inst.latch_mem_inst.gen_gclk\[44\]._gclk
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.gclk\[44\] sky130_fd_sc_hd__clkbuf_4
X_2310_ net358 _0969_ _0977_ VGND VGND VDPWR VDPWR _0070_ sky130_fd_sc_hd__mux2_1
X_2172_ _0768_ _0817_ net167 VGND VGND VDPWR VDPWR _0862_ sky130_fd_sc_hd__o21a_1
X_2241_ _0230_ _0927_ VGND VGND VDPWR VDPWR _0928_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_48_453 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1956_ dig_ctrl_inst.latch_mem_inst.RAM\[46\]\[6\] net73 net57 _0145_ dig_ctrl_inst.latch_mem_inst.RAM\[45\]\[6\]
+ VGND VGND VDPWR VDPWR _0662_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_31_353 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[57\].gen_latches\[4\].p_latch net210 dig_ctrl_inst.latch_mem_inst.gclk\[57\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[57\]\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_7_113 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_1887_ dig_ctrl_inst.latch_mem_inst.RAM\[13\]\[5\] _0114_ _0150_ dig_ctrl_inst.latch_mem_inst.RAM\[52\]\[5\]
+ VGND VGND VDPWR VDPWR _0594_ sky130_fd_sc_hd__a22o_1
X_2508_ clknet_leaf_5_clk _0105_ net178 VGND VGND VDPWR VDPWR net19 sky130_fd_sc_hd__dfrtp_1
Xoutput19 net19 VGND VGND VDPWR VDPWR port_ms_o[2] sky130_fd_sc_hd__buf_2
XFILLER_0_3_341 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_2439_ clknet_leaf_8_clk _0047_ net146 VGND VGND VDPWR VDPWR dig_ctrl_inst.cpu_inst.r0\[2\]
+ sky130_fd_sc_hd__dfrtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[46\].gen_latches\[2\].p_latch net228 dig_ctrl_inst.latch_mem_inst.gclk\[46\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[46\]\[2\] sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_54_489 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2527__274 VGND VGND VDPWR VDPWR _2527__274/HI net274 sky130_fd_sc_hd__conb_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[1\].gen_latches\[6\].p_latch net195 dig_ctrl_inst.latch_mem_inst.gclk\[1\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[1\]\[6\] sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[35\].gen_latches\[0\].p_latch net240 dig_ctrl_inst.latch_mem_inst.gclk\[35\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[35\]\[0\] sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_45_434 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_15 VDPWR VGND VDPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_306 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
X_1741_ dig_ctrl_inst.latch_mem_inst.RAM\[44\]\[3\] _0144_ _0146_ dig_ctrl_inst.latch_mem_inst.RAM\[47\]\[3\]
+ VGND VGND VDPWR VDPWR _0450_ sky130_fd_sc_hd__a22o_1
X_1810_ _0512_ _0513_ _0517_ VGND VGND VDPWR VDPWR _0518_ sky130_fd_sc_hd__or3_1
X_1672_ dig_ctrl_inst.latch_mem_inst.RAM\[11\]\[1\] _1145_ _0126_ dig_ctrl_inst.latch_mem_inst.RAM\[23\]\[1\]
+ _0377_ VGND VGND VDPWR VDPWR _0383_ sky130_fd_sc_hd__a221o_1
XFILLER_0_40_203 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_333 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[23\].gen_latches\[7\].p_latch net183 dig_ctrl_inst.latch_mem_inst.gclk\[23\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[23\]\[7\] sky130_fd_sc_hd__dlxtp_1
X_2224_ net160 _0890_ VGND VGND VDPWR VDPWR _0912_ sky130_fd_sc_hd__xnor2_1
X_2155_ net168 _0786_ _0783_ net169 VGND VGND VDPWR VDPWR _0846_ sky130_fd_sc_hd__a2bb2o_1
X_2086_ _0233_ net137 VGND VGND VDPWR VDPWR _0779_ sky130_fd_sc_hd__nand2_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[12\].gen_latches\[5\].p_latch net200 dig_ctrl_inst.latch_mem_inst.gclk\[12\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[12\]\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_31_247 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_225 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
X_1939_ dig_ctrl_inst.latch_mem_inst.RAM\[26\]\[6\] net84 net65 VGND VGND VDPWR VDPWR
+ _0645_ sky130_fd_sc_hd__and3_2
XFILLER_0_16_244 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_8
Xdig_ctrl_inst.latch_mem_inst.gen_words\[5\].gen_latches\[7\].p_latch net187 dig_ctrl_inst.latch_mem_inst.gclk\[5\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[5\]\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_66_133 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_415 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_11_Right_11 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[39\].gen_latches\[1\].p_latch net232 dig_ctrl_inst.latch_mem_inst.gclk\[39\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[39\]\[1\] sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[1\].clock_buffer dig_ctrl_inst.latch_mem_inst.gen_gclk\[1\]._gclk
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.gclk\[1\] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_38_26 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_20_Right_20 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_111 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
Xhold104 net20 VGND VGND VDPWR VDPWR net386 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_309 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
X_1724_ _0417_ _0419_ _0423_ _0433_ VGND VGND VDPWR VDPWR _0434_ sky130_fd_sc_hd__or4_1
X_1586_ dig_ctrl_inst.latch_mem_inst.RAM\[10\]\[0\] net121 net294 VGND VGND VDPWR
+ VDPWR _0298_ sky130_fd_sc_hd__and3_2
X_1655_ dig_ctrl_inst.latch_mem_inst.RAM\[16\]\[1\] net128 net61 VGND VGND VDPWR VDPWR
+ _0366_ sky130_fd_sc_hd__and3_2
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[17\].clock_gate clknet_leaf_1_clk dig_ctrl_inst.latch_mem_inst.data_we\[17\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.gen_gclk\[17\]._gclk sky130_fd_sc_hd__dlclkp_1
XTAP_TAPCELL_ROW_64_551 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_111 VDPWR VGND VDPWR VGND sky130_ef_sc_hd__decap_12
X_2138_ _0828_ _0829_ VGND VGND VDPWR VDPWR _0830_ sky130_fd_sc_hd__and2_1
XFILLER_0_28_81 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
X_2069_ net166 net137 VGND VGND VDPWR VDPWR _0762_ sky130_fd_sc_hd__nand2_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[16\].gen_latches\[6\].p_latch net191 dig_ctrl_inst.latch_mem_inst.gclk\[16\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[16\]\[6\] sky130_fd_sc_hd__dlxtp_1
X_2207_ _1118_ _0790_ _0825_ net169 VGND VGND VDPWR VDPWR _0896_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_21_3 VDPWR VGND VDPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_169 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_125 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_166 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_111 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_70_587 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1371_ net83 net60 VGND VGND VDPWR VDPWR _0142_ sky130_fd_sc_hd__and2_2
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[37\].clock_buffer dig_ctrl_inst.latch_mem_inst.gen_gclk\[37\]._gclk
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.gclk\[37\] sky130_fd_sc_hd__clkbuf_4
X_1440_ net248 _1007_ dig_ctrl_inst.cpu_inst.prev_state\[2\] _0999_ VGND VGND VDPWR
+ VDPWR _0177_ sky130_fd_sc_hd__a22o_1
XFILLER_0_4_27 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_532 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_136 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_317 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_275 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_3 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
X_1707_ dig_ctrl_inst.latch_mem_inst.RAM\[24\]\[2\] _0127_ _0136_ dig_ctrl_inst.latch_mem_inst.RAM\[34\]\[2\]
+ VGND VGND VDPWR VDPWR _0417_ sky130_fd_sc_hd__a22o_1
X_1638_ dig_ctrl_inst.latch_mem_inst.RAM\[18\]\[1\] net109 net61 VGND VGND VDPWR VDPWR
+ _0349_ sky130_fd_sc_hd__and3_2
X_1569_ _1048_ net108 net123 VGND VGND VDPWR VDPWR _0281_ sky130_fd_sc_hd__a21bo_1
XPHY_EDGE_ROW_18_Left_96 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
Xfanout98 _1137_ VGND VGND VDPWR VDPWR net98 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_44_180 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
Xfanout87 _1141_ VGND VGND VDPWR VDPWR net87 sky130_fd_sc_hd__buf_2
Xfanout65 net66 VGND VGND VDPWR VDPWR net65 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout54 net60 VGND VGND VDPWR VDPWR net54 sky130_fd_sc_hd__buf_6
Xfanout76 net79 VGND VGND VDPWR VDPWR net76 sky130_fd_sc_hd__clkbuf_2
Xfanout43 net44 VGND VGND VDPWR VDPWR net43 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_9_221 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_17 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_75_613 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_169 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_125 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_15_256 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2472_ clknet_leaf_4_clk _0078_ VGND VGND VDPWR VDPWR dig_ctrl_inst.spi_receiver_inst.stb_o
+ sky130_fd_sc_hd__dfxtp_1
Xclkload13 clknet_leaf_6_clk VGND VGND VDPWR VDPWR clkload13/Y sky130_fd_sc_hd__clkinv_8
XFILLER_0_35_180 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_9 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_1285_ net304 _1078_ net301 VGND VGND VDPWR VDPWR _1131_ sky130_fd_sc_hd__a21oi_1
X_1423_ net255 dig_ctrl_inst.cpu_inst.r1\[6\] VGND VGND VDPWR VDPWR _0165_ sky130_fd_sc_hd__and2b_1
X_1354_ net128 net150 net55 VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.data_we\[32\]
+ sky130_fd_sc_hd__and3_2
Xclkload7 clknet_leaf_18_clk VGND VGND VDPWR VDPWR clkload7/Y sky130_fd_sc_hd__inv_16
XFILLER_0_14_331 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_114 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
Xfanout222 net223 VGND VGND VDPWR VDPWR net222 sky130_fd_sc_hd__buf_2
Xfanout211 net213 VGND VGND VDPWR VDPWR net211 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_41_172 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_8
Xfanout200 net201 VGND VGND VDPWR VDPWR net200 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_TAPCELL_ROW_6_202 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout244 net245 VGND VGND VDPWR VDPWR net244 sky130_fd_sc_hd__clkbuf_2
Xfanout255 dig_ctrl_inst.cpu_inst.arg1\[1\] VGND VGND VDPWR VDPWR net255 sky130_fd_sc_hd__clkbuf_2
Xfanout266 dig_ctrl_inst.cpu_inst.arg0\[0\] VGND VGND VDPWR VDPWR net266 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_29_337 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout233 net327 VGND VGND VDPWR VDPWR net233 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_12_237 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_59 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_26 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_39 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
X_1972_ dig_ctrl_inst.latch_mem_inst.RAM\[15\]\[6\] _0117_ _0625_ _0636_ _0658_ VGND
+ VGND VDPWR VDPWR _0678_ sky130_fd_sc_hd__a2111o_1
X_2524_ net273 VGND VGND VDPWR VDPWR uio_oe[5] sky130_fd_sc_hd__buf_2
XFILLER_0_70_256 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_49_Right_49 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
X_2455_ clknet_leaf_8_clk _0063_ net143 VGND VGND VDPWR VDPWR dig_ctrl_inst.cpu_inst.r2\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_11_73 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_312 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_2386_ clknet_leaf_3_clk net6 net174 VGND VGND VDPWR VDPWR dig_ctrl_inst.synchronizer_port_i_inst\[3\].pipe\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_58_Right_58 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
X_1268_ net256 dig_ctrl_inst.cpu_inst.r1\[4\] VGND VGND VDPWR VDPWR _1116_ sky130_fd_sc_hd__and2b_1
X_1406_ net115 net80 net44 VGND VGND VDPWR VDPWR _0158_ sky130_fd_sc_hd__and3_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[53\].gen_latches\[7\].p_latch net184 dig_ctrl_inst.latch_mem_inst.gclk\[53\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[53\]\[7\] sky130_fd_sc_hd__dlxtp_1
X_1337_ net150 _0126_ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.data_we\[23\]
+ sky130_fd_sc_hd__and2_1
X_1199_ net249 _1029_ _1038_ _1046_ _1008_ VGND VGND VDPWR VDPWR _1047_ sky130_fd_sc_hd__o41a_4
XTAP_TAPCELL_ROW_26_318 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_67_Right_67 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[42\].gen_latches\[5\].p_latch net205 dig_ctrl_inst.latch_mem_inst.gclk\[42\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[42\]\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_14_172 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_76_Right_76 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[31\].gen_latches\[3\].p_latch net215 dig_ctrl_inst.latch_mem_inst.gclk\[31\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[31\]\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_37_275 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[20\].gen_latches\[1\].p_latch net235 dig_ctrl_inst.latch_mem_inst.gclk\[20\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[20\]\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_20_120 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
X_2171_ _0768_ _0808_ _0816_ _0765_ VGND VGND VDPWR VDPWR _0861_ sky130_fd_sc_hd__o22a_1
X_2240_ _0244_ _0906_ _0241_ VGND VGND VDPWR VDPWR _0927_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_75_337 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_48_454 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_103 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
X_1955_ dig_ctrl_inst.latch_mem_inst.RAM\[21\]\[6\] _0124_ _0277_ dig_ctrl_inst.latch_mem_inst.RAM\[4\]\[6\]
+ VGND VGND VDPWR VDPWR _0661_ sky130_fd_sc_hd__a22o_1
X_1886_ _0582_ _0586_ _0588_ _0592_ VGND VGND VDPWR VDPWR _0593_ sky130_fd_sc_hd__or4_1
XFILLER_0_7_147 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
X_2507_ clknet_leaf_4_clk _0104_ net178 VGND VGND VDPWR VDPWR net18 sky130_fd_sc_hd__dfrtp_1
X_2438_ clknet_leaf_7_clk _0046_ net144 VGND VGND VDPWR VDPWR dig_ctrl_inst.cpu_inst.r0\[1\]
+ sky130_fd_sc_hd__dfrtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[2\].gen_latches\[1\].p_latch net232 dig_ctrl_inst.latch_mem_inst.gclk\[2\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[2\]\[1\] sky130_fd_sc_hd__dlxtp_1
X_2369_ net253 _1013_ _0175_ net252 VGND VGND VDPWR VDPWR _0996_ sky130_fd_sc_hd__and4b_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[46\].gen_latches\[6\].p_latch net197 dig_ctrl_inst.latch_mem_inst.gclk\[46\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[46\]\[6\] sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[35\].gen_latches\[4\].p_latch net210 dig_ctrl_inst.latch_mem_inst.gclk\[35\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[35\]\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_6_191 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[24\].clock_gate clknet_leaf_17_clk dig_ctrl_inst.latch_mem_inst.data_we\[24\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.gen_gclk\[24\]._gclk sky130_fd_sc_hd__dlclkp_1
XFILLER_0_27_17 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_337 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_45_435 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_49 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_27 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[24\].gen_latches\[2\].p_latch net227 dig_ctrl_inst.latch_mem_inst.gclk\[24\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[24\]\[2\] sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_6_Left_84 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
X_1671_ dig_ctrl_inst.latch_mem_inst.RAM\[3\]\[1\] _1135_ _0130_ dig_ctrl_inst.latch_mem_inst.RAM\[27\]\[1\]
+ _0378_ VGND VGND VDPWR VDPWR _0382_ sky130_fd_sc_hd__a221o_1
X_1740_ net261 _0449_ _0276_ VGND VGND VDPWR VDPWR _0028_ sky130_fd_sc_hd__mux2_1
XFILLER_0_25_223 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_24 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[13\].gen_latches\[0\].p_latch net246 dig_ctrl_inst.latch_mem_inst.gclk\[13\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[13\]\[0\] sky130_fd_sc_hd__dlxtp_1
X_2223_ net160 net159 _0867_ VGND VGND VDPWR VDPWR _0911_ sky130_fd_sc_hd__or3_1
X_2154_ _0748_ _0750_ _0844_ VGND VGND VDPWR VDPWR _0845_ sky130_fd_sc_hd__mux2_1
X_2085_ net138 net137 net157 VGND VGND VDPWR VDPWR _0778_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_17_61 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_223 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_8
X_1938_ dig_ctrl_inst.latch_mem_inst.RAM\[56\]\[6\] net88 net48 VGND VGND VDPWR VDPWR
+ _0644_ sky130_fd_sc_hd__and3_2
X_1869_ dig_ctrl_inst.latch_mem_inst.RAM\[29\]\[5\] _0131_ _0277_ dig_ctrl_inst.latch_mem_inst.RAM\[4\]\[5\]
+ VGND VGND VDPWR VDPWR _0576_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_59_516 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[6\].gen_latches\[2\].p_latch net226 dig_ctrl_inst.latch_mem_inst.gclk\[6\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[6\]\[2\] sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_42_416 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_337 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[39\].gen_latches\[5\].p_latch net206 dig_ctrl_inst.latch_mem_inst.gclk\[39\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[39\]\[5\] sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[28\].gen_latches\[3\].p_latch net222 dig_ctrl_inst.latch_mem_inst.gclk\[28\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[28\]\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_54_59 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_126 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_318 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
X_1723_ dig_ctrl_inst.latch_mem_inst.RAM\[36\]\[2\] net96 net58 _0279_ dig_ctrl_inst.latch_mem_inst.RAM\[6\]\[2\]
+ VGND VGND VDPWR VDPWR _0433_ sky130_fd_sc_hd__a32o_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[17\].gen_latches\[1\].p_latch net239 dig_ctrl_inst.latch_mem_inst.gclk\[17\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[17\]\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_13_248 VDPWR VGND VDPWR VGND sky130_ef_sc_hd__decap_12
Xhold105 dig_ctrl_inst.cpu_inst.data\[7\] VGND VGND VDPWR VDPWR net387 sky130_fd_sc_hd__dlygate4sd3_1
X_1654_ dig_ctrl_inst.latch_mem_inst.RAM\[10\]\[1\] net121 net294 VGND VGND VDPWR
+ VDPWR _0365_ sky130_fd_sc_hd__and3_2
XFILLER_0_0_197 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_2206_ _0238_ _0792_ _0894_ VGND VGND VDPWR VDPWR _0895_ sky130_fd_sc_hd__a21oi_1
X_1585_ dig_ctrl_inst.latch_mem_inst.RAM\[25\]\[0\] net116 net90 net63 VGND VGND VDPWR
+ VDPWR _0297_ sky130_fd_sc_hd__and4_1
X_2137_ net165 net162 VGND VGND VDPWR VDPWR _0829_ sky130_fd_sc_hd__nand2_1
XFILLER_0_44_81 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
X_2068_ net169 net137 VGND VGND VDPWR VDPWR _0761_ sky130_fd_sc_hd__nand2_1
XFILLER_0_14_3 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_220 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_189 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_29 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_15 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_48 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_8
X_1370_ net152 _0141_ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.data_we\[41\]
+ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_61_533 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_126 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_62 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_307 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_1706_ dig_ctrl_inst.latch_mem_inst.RAM\[7\]\[2\] net126 net106 net101 VGND VGND
+ VDPWR VDPWR _0416_ sky130_fd_sc_hd__and4_1
XFILLER_0_5_256 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_6
X_1637_ dig_ctrl_inst.latch_mem_inst.RAM\[38\]\[1\] net94 net54 VGND VGND VDPWR VDPWR
+ _0348_ sky130_fd_sc_hd__and3_2
X_1568_ net119 _1131_ net101 net123 VGND VGND VDPWR VDPWR _0280_ sky130_fd_sc_hd__o211a_1
X_1499_ dig_ctrl_inst.cpu_inst.ip\[0\] dig_ctrl_inst.cpu_inst.ip\[1\] dig_ctrl_inst.cpu_inst.ip\[2\]
+ dig_ctrl_inst.cpu_inst.ip\[3\] VGND VGND VDPWR VDPWR _0215_ sky130_fd_sc_hd__and4_1
Xfanout55 net60 VGND VGND VDPWR VDPWR net55 sky130_fd_sc_hd__clkbuf_2
Xfanout44 net47 VGND VGND VDPWR VDPWR net44 sky130_fd_sc_hd__buf_2
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[3\].clock_gate clknet_leaf_3_clk dig_ctrl_inst.latch_mem_inst.data_we\[3\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.gen_gclk\[3\]._gclk sky130_fd_sc_hd__dlclkp_1
Xfanout88 net89 VGND VGND VDPWR VDPWR net88 sky130_fd_sc_hd__buf_2
Xfanout77 net79 VGND VGND VDPWR VDPWR net77 sky130_fd_sc_hd__buf_1
Xfanout66 net67 VGND VGND VDPWR VDPWR net66 sky130_fd_sc_hd__buf_4
Xfanout99 net100 VGND VGND VDPWR VDPWR net99 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_3_3 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_75_614 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[61\].gen_latches\[3\].p_latch net215 dig_ctrl_inst.latch_mem_inst.gclk\[61\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[61\]\[3\] sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_15_257 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2471_ clknet_leaf_3_clk _0077_ net173 VGND VGND VDPWR VDPWR dig_ctrl_inst.spi_miso_o
+ sky130_fd_sc_hd__dfrtp_1
Xclkload14 clknet_leaf_7_clk VGND VGND VDPWR VDPWR clkload14/Y sky130_fd_sc_hd__clkinv_16
X_1422_ net259 dig_ctrl_inst.cpu_inst.r2\[6\] VGND VGND VDPWR VDPWR _0164_ sky130_fd_sc_hd__and2b_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[50\].gen_latches\[1\].p_latch net232 dig_ctrl_inst.latch_mem_inst.gclk\[50\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[50\]\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_23_332 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
XFILLER_0_76_57 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_1284_ net154 _1130_ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.data_we\[1\]
+ sky130_fd_sc_hd__and2_1
X_1353_ net129 net53 VGND VGND VDPWR VDPWR _0134_ sky130_fd_sc_hd__and2_2
XFILLER_0_58_273 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
Xclkload8 clknet_leaf_1_clk VGND VGND VDPWR VDPWR clkload8/Y sky130_fd_sc_hd__inv_12
XFILLER_0_41_71 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[29\].clock_gate clknet_leaf_0_clk dig_ctrl_inst.latch_mem_inst.data_we\[29\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.gen_gclk\[29\]._gclk sky130_fd_sc_hd__dlclkp_1
Xfanout245 net246 VGND VGND VDPWR VDPWR net245 sky130_fd_sc_hd__clkbuf_2
Xfanout223 net329 VGND VGND VDPWR VDPWR net223 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout212 net213 VGND VGND VDPWR VDPWR net212 sky130_fd_sc_hd__clkbuf_2
Xfanout256 net257 VGND VGND VDPWR VDPWR net256 sky130_fd_sc_hd__buf_4
Xfanout234 net236 VGND VGND VDPWR VDPWR net234 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_1_281 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_6_203 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout201 net202 VGND VGND VDPWR VDPWR net201 sky130_fd_sc_hd__clkbuf_2
Xfanout267 net268 VGND VGND VDPWR VDPWR net267 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_29_338 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_238 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_282 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[31\].clock_gate clknet_leaf_15_clk dig_ctrl_inst.latch_mem_inst.data_we\[31\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.gen_gclk\[31\]._gclk sky130_fd_sc_hd__dlclkp_1
X_1971_ dig_ctrl_inst.latch_mem_inst.RAM\[13\]\[6\] _0114_ _0630_ _0641_ _0657_ VGND
+ VGND VDPWR VDPWR _0677_ sky130_fd_sc_hd__a2111o_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[54\].gen_latches\[2\].p_latch net224 dig_ctrl_inst.latch_mem_inst.gclk\[54\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[54\]\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_23_140 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
X_2523_ net272 VGND VGND VDPWR VDPWR uio_oe[4] sky130_fd_sc_hd__buf_2
X_2520__270 VGND VGND VDPWR VDPWR _2520__270/HI net270 sky130_fd_sc_hd__conb_1
X_1405_ net153 net78 net48 VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.data_we\[60\]
+ sky130_fd_sc_hd__and3_2
X_2385_ clknet_leaf_4_clk net332 net174 VGND VGND VDPWR VDPWR dig_ctrl_inst.synchronizer_port_i_inst\[4\].out
+ sky130_fd_sc_hd__dfrtp_1
X_2454_ clknet_leaf_9_clk _0062_ net141 VGND VGND VDPWR VDPWR dig_ctrl_inst.cpu_inst.r2\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_11_335 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_1198_ _1039_ _1045_ VGND VGND VDPWR VDPWR _1046_ sky130_fd_sc_hd__and2_1
X_1267_ net260 net256 dig_ctrl_inst.cpu_inst.r2\[4\] VGND VGND VDPWR VDPWR _1115_
+ sky130_fd_sc_hd__and3b_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[43\].gen_latches\[0\].p_latch net245 dig_ctrl_inst.latch_mem_inst.gclk\[43\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[43\]\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_36_82 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_71 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_26_319 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1336_ net102 net99 net63 VGND VGND VDPWR VDPWR _0126_ sky130_fd_sc_hd__and3_4
Xinput1 port_ms_i VGND VGND VDPWR VDPWR net1 sky130_fd_sc_hd__buf_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[31\].gen_latches\[7\].p_latch net187 dig_ctrl_inst.latch_mem_inst.gclk\[31\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[31\]\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_32_29 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_257 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[20\].gen_latches\[5\].p_latch net207 dig_ctrl_inst.latch_mem_inst.gclk\[20\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[20\]\[5\] sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_48_455 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2170_ _0809_ _0836_ _0859_ _0770_ VGND VGND VDPWR VDPWR _0860_ sky130_fd_sc_hd__o22a_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[58\].gen_latches\[3\].p_latch net223 dig_ctrl_inst.latch_mem_inst.gclk\[58\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[58\]\[3\] sky130_fd_sc_hd__dlxtp_1
X_1954_ dig_ctrl_inst.latch_mem_inst.RAM\[22\]\[6\] _0125_ _0153_ dig_ctrl_inst.latch_mem_inst.RAM\[55\]\[6\]
+ VGND VGND VDPWR VDPWR _0660_ sky130_fd_sc_hd__a22o_1
XFILLER_0_43_202 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_1885_ dig_ctrl_inst.latch_mem_inst.RAM\[3\]\[5\] _1135_ _0589_ _0590_ _0591_ VGND
+ VGND VDPWR VDPWR _0592_ sky130_fd_sc_hd__a2111o_1
X_2506_ clknet_leaf_3_clk _0103_ net178 VGND VGND VDPWR VDPWR net17 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_44_3 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_2437_ clknet_leaf_7_clk _0045_ net144 VGND VGND VDPWR VDPWR dig_ctrl_inst.cpu_inst.r0\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_39_400 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2368_ _0566_ _0991_ _0992_ _0993_ _0994_ VGND VGND VDPWR VDPWR _0995_ sky130_fd_sc_hd__a2111o_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[47\].gen_latches\[1\].p_latch net236 dig_ctrl_inst.latch_mem_inst.gclk\[47\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[47\]\[1\] sky130_fd_sc_hd__dlxtp_1
X_1319_ net126 net106 net82 VGND VGND VDPWR VDPWR _0117_ sky130_fd_sc_hd__and3_4
X_2299_ _1024_ _0175_ _0756_ VGND VGND VDPWR VDPWR _0976_ sky130_fd_sc_hd__and3_4
XFILLER_0_2_83 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[2\].gen_latches\[5\].p_latch net203 dig_ctrl_inst.latch_mem_inst.gclk\[2\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[2\]\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_34_213 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_181 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XFILLER_0_69_121 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
Xmax_cap85 _1144_ VGND VGND VDPWR VDPWR net85 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_TAPCELL_ROW_53_480 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_436 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[24\].gen_latches\[6\].p_latch net194 dig_ctrl_inst.latch_mem_inst.gclk\[24\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[24\]\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_4_118 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_28 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
X_1670_ dig_ctrl_inst.latch_mem_inst.RAM\[55\]\[1\] _0153_ _0341_ _0359_ _0360_ VGND
+ VGND VDPWR VDPWR _0381_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_68_36 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
X_2222_ net167 _0810_ _0819_ _0909_ net171 VGND VGND VDPWR VDPWR _0910_ sky130_fd_sc_hd__a221o_1
XFILLER_0_48_316 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[13\].gen_latches\[4\].p_latch net211 dig_ctrl_inst.latch_mem_inst.gclk\[13\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[13\]\[4\] sky130_fd_sc_hd__dlxtp_1
X_2084_ _0775_ _0776_ _1068_ VGND VGND VDPWR VDPWR _0777_ sky130_fd_sc_hd__mux2_1
X_2153_ _0842_ _0843_ VGND VGND VDPWR VDPWR _0844_ sky130_fd_sc_hd__nand2_1
X_1937_ dig_ctrl_inst.latch_mem_inst.RAM\[34\]\[6\] net110 net55 VGND VGND VDPWR VDPWR
+ _0643_ sky130_fd_sc_hd__and3_2
XFILLER_0_16_257 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[40\].clock_buffer dig_ctrl_inst.latch_mem_inst.gen_gclk\[40\]._gclk
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.gclk\[40\] sky130_fd_sc_hd__clkbuf_4
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[8\].clock_gate clknet_leaf_3_clk dig_ctrl_inst.latch_mem_inst.data_we\[8\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.gen_gclk\[8\]._gclk sky130_fd_sc_hd__dlclkp_1
X_1868_ dig_ctrl_inst.latch_mem_inst.RAM\[59\]\[5\] _0156_ _0279_ dig_ctrl_inst.latch_mem_inst.RAM\[6\]\[5\]
+ VGND VGND VDPWR VDPWR _0575_ sky130_fd_sc_hd__a22o_1
X_1799_ dig_ctrl_inst.latch_mem_inst.RAM\[17\]\[4\] _0120_ _0127_ dig_ctrl_inst.latch_mem_inst.RAM\[24\]\[4\]
+ VGND VGND VDPWR VDPWR _0507_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_59_517 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_417 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_327 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[6\].gen_latches\[6\].p_latch net194 dig_ctrl_inst.latch_mem_inst.gclk\[6\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[6\]\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_15_290 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_27 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[28\].gen_latches\[7\].p_latch net185 dig_ctrl_inst.latch_mem_inst.gclk\[28\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[28\]\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_70_26 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_341 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_1722_ dig_ctrl_inst.latch_mem_inst.RAM\[51\]\[2\] _0149_ _0277_ dig_ctrl_inst.latch_mem_inst.RAM\[4\]\[2\]
+ _0402_ VGND VGND VDPWR VDPWR _0432_ sky130_fd_sc_hd__a221o_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[17\].gen_latches\[5\].p_latch net202 dig_ctrl_inst.latch_mem_inst.gclk\[17\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[17\]\[5\] sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_9_Right_9 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
X_1584_ dig_ctrl_inst.latch_mem_inst.RAM\[28\]\[0\] net76 net63 VGND VGND VDPWR VDPWR
+ _0296_ sky130_fd_sc_hd__and3_2
Xhold106 dig_ctrl_inst.cpu_inst.data\[6\] VGND VGND VDPWR VDPWR net388 sky130_fd_sc_hd__dlygate4sd3_1
X_1653_ dig_ctrl_inst.latch_mem_inst.RAM\[36\]\[1\] net96 net56 VGND VGND VDPWR VDPWR
+ _0364_ sky130_fd_sc_hd__and3_2
XFILLER_0_0_187 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_2205_ dig_ctrl_inst.cpu_inst.data\[4\] _0743_ _0783_ net160 VGND VGND VDPWR VDPWR
+ _0894_ sky130_fd_sc_hd__a22o_1
XFILLER_0_48_168 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_135 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
X_2136_ net165 net162 VGND VGND VDPWR VDPWR _0828_ sky130_fd_sc_hd__or2_1
XFILLER_0_8_210 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
X_2067_ _1103_ _1118_ _0167_ _0172_ VGND VGND VDPWR VDPWR _0760_ sky130_fd_sc_hd__or4_2
XPHY_EDGE_ROW_22_Left_100 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_4_186 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[36\].clock_gate clknet_leaf_19_clk dig_ctrl_inst.latch_mem_inst.data_we\[36\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.gen_gclk\[36\]._gclk sky130_fd_sc_hd__dlclkp_1
XFILLER_0_54_138 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_113 VDPWR VGND VDPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_341 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_311 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_1705_ dig_ctrl_inst.latch_mem_inst.RAM\[44\]\[2\] net77 net54 VGND VGND VDPWR VDPWR
+ _0415_ sky130_fd_sc_hd__and3_2
XFILLER_0_5_279 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_74 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_1567_ net125 net95 VGND VGND VDPWR VDPWR _0279_ sky130_fd_sc_hd__and2_2
X_1636_ dig_ctrl_inst.latch_mem_inst.RAM\[48\]\[1\] net130 net46 VGND VGND VDPWR VDPWR
+ _0347_ sky130_fd_sc_hd__and3_2
X_1498_ _0214_ _0204_ dig_ctrl_inst.cpu_inst.ip\[2\] _0211_ VGND VGND VDPWR VDPWR
+ _0021_ sky130_fd_sc_hd__a2bb2o_1
X_2119_ _0762_ _0766_ _1068_ VGND VGND VDPWR VDPWR _0811_ sky130_fd_sc_hd__mux2_1
Xfanout78 net79 VGND VGND VDPWR VDPWR net78 sky130_fd_sc_hd__buf_2
Xfanout67 _0118_ VGND VGND VDPWR VDPWR net67 sky130_fd_sc_hd__buf_4
Xfanout56 net60 VGND VGND VDPWR VDPWR net56 sky130_fd_sc_hd__clkbuf_2
Xfanout45 net47 VGND VGND VDPWR VDPWR net45 sky130_fd_sc_hd__buf_2
XFILLER_0_44_160 VDPWR VGND VDPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_341 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_75_615 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload15 clknet_leaf_8_clk VGND VGND VDPWR VDPWR clkload15/Y sky130_fd_sc_hd__inv_12
Xdig_ctrl_inst.latch_mem_inst.gen_words\[61\].gen_latches\[7\].p_latch net184 dig_ctrl_inst.latch_mem_inst.gclk\[61\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[61\]\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_76_36 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
X_1421_ net259 net255 dig_ctrl_inst.cpu_inst.r3\[6\] VGND VGND VDPWR VDPWR _0163_
+ sky130_fd_sc_hd__and3_2
X_2470_ clknet_leaf_11_clk _0076_ net140 VGND VGND VDPWR VDPWR dig_ctrl_inst.cpu_inst.r3\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_1283_ net132 net125 net118 VGND VGND VDPWR VDPWR _1130_ sky130_fd_sc_hd__and3_2
X_1352_ _1127_ _1112_ VGND VGND VDPWR VDPWR _0133_ sky130_fd_sc_hd__and2b_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[50\].gen_latches\[5\].p_latch net203 dig_ctrl_inst.latch_mem_inst.gclk\[50\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[50\]\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_73_222 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_241 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[33\].clock_buffer dig_ctrl_inst.latch_mem_inst.gen_gclk\[33\]._gclk
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.gclk\[33\] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_74_3 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
Xclkload9 clknet_leaf_2_clk VGND VGND VDPWR VDPWR clkload9/Y sky130_fd_sc_hd__inv_16
Xfanout213 net214 VGND VGND VDPWR VDPWR net213 sky130_fd_sc_hd__buf_2
X_1619_ _0327_ _0328_ _0329_ _0330_ VGND VGND VDPWR VDPWR _0331_ sky130_fd_sc_hd__or4_1
Xfanout246 net247 VGND VGND VDPWR VDPWR net246 sky130_fd_sc_hd__buf_2
Xfanout268 dig_ctrl_inst.cpu_inst.arg0\[0\] VGND VGND VDPWR VDPWR net268 sky130_fd_sc_hd__buf_4
Xfanout257 dig_ctrl_inst.cpu_inst.arg1\[1\] VGND VGND VDPWR VDPWR net257 sky130_fd_sc_hd__buf_2
Xfanout202 net207 VGND VGND VDPWR VDPWR net202 sky130_fd_sc_hd__buf_2
Xfanout235 net236 VGND VGND VDPWR VDPWR net235 sky130_fd_sc_hd__buf_1
Xfanout224 net225 VGND VGND VDPWR VDPWR net224 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_29_339 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_239 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_283 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1970_ dig_ctrl_inst.latch_mem_inst.RAM\[31\]\[6\] _0132_ _0134_ dig_ctrl_inst.latch_mem_inst.RAM\[32\]\[6\]
+ _0643_ VGND VGND VDPWR VDPWR _0676_ sky130_fd_sc_hd__a221o_1
X_2522_ net271 VGND VGND VDPWR VDPWR uio_oe[3] sky130_fd_sc_hd__buf_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[54\].gen_latches\[6\].p_latch net191 dig_ctrl_inst.latch_mem_inst.gclk\[54\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[54\]\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_15_119 VDPWR VGND VDPWR VGND sky130_ef_sc_hd__decap_12
X_2384_ clknet_leaf_3_clk net7 net174 VGND VGND VDPWR VDPWR dig_ctrl_inst.synchronizer_port_i_inst\[4\].pipe\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_1404_ net78 net49 VGND VGND VDPWR VDPWR _0157_ sky130_fd_sc_hd__and2_2
X_1335_ net149 net93 net61 VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.data_we\[22\]
+ sky130_fd_sc_hd__and3_2
X_2453_ clknet_leaf_11_clk _0061_ net140 VGND VGND VDPWR VDPWR dig_ctrl_inst.cpu_inst.r2\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xinput2 rst_n VGND VGND VDPWR VDPWR net2 sky130_fd_sc_hd__clkbuf_1
X_1266_ net261 net256 dig_ctrl_inst.cpu_inst.r3\[4\] VGND VGND VDPWR VDPWR _1114_
+ sky130_fd_sc_hd__and3_2
X_1197_ net300 _1041_ _1042_ _1043_ _1044_ VGND VGND VDPWR VDPWR _1045_ sky130_fd_sc_hd__o41a_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[43\].gen_latches\[4\].p_latch net213 dig_ctrl_inst.latch_mem_inst.gclk\[43\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[43\]\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_6_341 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[32\].gen_latches\[2\].p_latch net224 dig_ctrl_inst.latch_mem_inst.gclk\[32\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[32\]\[2\] sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[21\].gen_latches\[0\].p_latch net246 dig_ctrl_inst.latch_mem_inst.gclk\[21\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[21\]\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_32_19 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_190 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_69_Left_147 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[58\].gen_latches\[7\].p_latch net188 dig_ctrl_inst.latch_mem_inst.gclk\[58\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[58\]\[7\] sky130_fd_sc_hd__dlxtp_1
X_1953_ dig_ctrl_inst.latch_mem_inst.RAM\[62\]\[6\] net73 net50 VGND VGND VDPWR VDPWR
+ _0659_ sky130_fd_sc_hd__and3_2
X_1884_ dig_ctrl_inst.latch_mem_inst.RAM\[48\]\[5\] net128 net44 VGND VGND VDPWR VDPWR
+ _0591_ sky130_fd_sc_hd__and3_2
XFILLER_0_22_85 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
X_2505_ clknet_leaf_5_clk _0102_ net178 VGND VGND VDPWR VDPWR net35 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_43_247 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_333 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[3\].gen_latches\[0\].p_latch net243 dig_ctrl_inst.latch_mem_inst.gclk\[3\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[3\]\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_47_93 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_6
X_2436_ clknet_leaf_9_clk _0044_ VGND VGND VDPWR VDPWR dig_ctrl_inst.cpu_inst.prev_state\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_39_401 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_3 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_2367_ _0449_ _0623_ VGND VGND VDPWR VDPWR _0994_ sky130_fd_sc_hd__and2_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[47\].gen_latches\[5\].p_latch net203 dig_ctrl_inst.latch_mem_inst.gclk\[47\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[47\]\[5\] sky130_fd_sc_hd__dlxtp_1
X_1318_ net148 net120 net72 VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.data_we\[14\]
+ sky130_fd_sc_hd__and3_2
X_2298_ net377 _0975_ _0967_ VGND VGND VDPWR VDPWR _0060_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_339 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
X_1249_ _1040_ _1096_ VGND VGND VDPWR VDPWR _1097_ sky130_fd_sc_hd__nand2_1
XFILLER_0_2_51 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[36\].gen_latches\[3\].p_latch net218 dig_ctrl_inst.latch_mem_inst.gclk\[36\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[36\]\[3\] sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_input_latches\[1\].n_latch dig_ctrl_inst.data_out\[1\]
+ clknet_leaf_2_clk VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.wdata\[1\]
+ sky130_fd_sc_hd__dlxtn_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[25\].gen_latches\[1\].p_latch net232 dig_ctrl_inst.latch_mem_inst.gclk\[25\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[25\]\[1\] sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_53_481 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_437 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_225 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_214 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_15 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[26\].clock_buffer dig_ctrl_inst.latch_mem_inst.gen_gclk\[26\]._gclk
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.gclk\[26\] sky130_fd_sc_hd__clkbuf_4
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[43\].clock_gate clknet_1_1__leaf_clk dig_ctrl_inst.latch_mem_inst.data_we\[43\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.gen_gclk\[43\]._gclk sky130_fd_sc_hd__dlclkp_1
X_2221_ _0836_ _0859_ _0908_ _0770_ _0886_ VGND VGND VDPWR VDPWR _0909_ sky130_fd_sc_hd__o221a_1
X_2152_ net164 net161 net166 VGND VGND VDPWR VDPWR _0843_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_48_306 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
X_2083_ net159 net137 VGND VGND VDPWR VDPWR _0776_ sky130_fd_sc_hd__nand2_1
X_1867_ dig_ctrl_inst.latch_mem_inst.RAM\[8\]\[5\] _1142_ _0571_ _0572_ _0573_ VGND
+ VGND VDPWR VDPWR _0574_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_63_309 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
X_1936_ dig_ctrl_inst.latch_mem_inst.RAM\[6\]\[6\] net121 net94 VGND VGND VDPWR VDPWR
+ _0642_ sky130_fd_sc_hd__and3_2
XFILLER_0_16_203 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_1798_ net257 _0505_ _0276_ VGND VGND VDPWR VDPWR _0029_ sky130_fd_sc_hd__mux2_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[7\].gen_latches\[1\].p_latch net239 dig_ctrl_inst.latch_mem_inst.gclk\[7\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[7\]\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_3_152 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_130 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_59_518 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2419_ clknet_leaf_8_clk _0027_ net143 VGND VGND VDPWR VDPWR dig_ctrl_inst.cpu_inst.arg0\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_42_418 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_306 VDPWR VGND VDPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_50_462 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[29\].gen_latches\[2\].p_latch net229 dig_ctrl_inst.latch_mem_inst.gclk\[29\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[29\]\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_38_29 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[18\].gen_latches\[0\].p_latch net242 dig_ctrl_inst.latch_mem_inst.gclk\[18\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[18\]\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_57_169 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
X_1721_ dig_ctrl_inst.latch_mem_inst.RAM\[40\]\[2\] _0140_ _0153_ dig_ctrl_inst.latch_mem_inst.RAM\[55\]\[2\]
+ _0430_ VGND VGND VDPWR VDPWR _0431_ sky130_fd_sc_hd__a221o_1
Xhold107 net29 VGND VGND VDPWR VDPWR net389 sky130_fd_sc_hd__dlygate4sd3_1
X_1583_ dig_ctrl_inst.latch_mem_inst.RAM\[27\]\[0\] net104 net91 net66 VGND VGND VDPWR
+ VDPWR _0295_ sky130_fd_sc_hd__and4_1
X_1652_ dig_ctrl_inst.latch_mem_inst.RAM\[6\]\[1\] net120 net93 VGND VGND VDPWR VDPWR
+ _0363_ sky130_fd_sc_hd__and3_2
XFILLER_0_0_111 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_2204_ _0747_ _0892_ VGND VGND VDPWR VDPWR _0893_ sky130_fd_sc_hd__nand2_1
X_2135_ net166 _0783_ _0826_ VGND VGND VDPWR VDPWR _0827_ sky130_fd_sc_hd__a21oi_1
X_2066_ _1103_ _1118_ _0167_ _0172_ VGND VGND VDPWR VDPWR _0759_ sky130_fd_sc_hd__nor4_1
X_1919_ dig_ctrl_inst.latch_mem_inst.RAM\[54\]\[6\] net93 net44 VGND VGND VDPWR VDPWR
+ _0625_ sky130_fd_sc_hd__and3_2
XFILLER_0_8_83 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_272 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_125 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_4_187 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1704_ dig_ctrl_inst.latch_mem_inst.RAM\[29\]\[2\] net119 _1146_ net69 VGND VGND
+ VDPWR VDPWR _0414_ sky130_fd_sc_hd__and4_1
XFILLER_0_60_109 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_85 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_214 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
X_1566_ net125 net118 net101 VGND VGND VDPWR VDPWR _0278_ sky130_fd_sc_hd__and3_2
XFILLER_0_39_72 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_1497_ _0173_ _0213_ _0212_ VGND VGND VDPWR VDPWR _0214_ sky130_fd_sc_hd__a21oi_1
X_1635_ dig_ctrl_inst.latch_mem_inst.RAM\[34\]\[1\] net109 net55 VGND VGND VDPWR VDPWR
+ _0346_ sky130_fd_sc_hd__and3_2
XTAP_TAPCELL_ROW_1_168 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2118_ _0770_ _0809_ VGND VGND VDPWR VDPWR _0810_ sky130_fd_sc_hd__or2_1
X_2049_ net252 net253 VGND VGND VDPWR VDPWR _0742_ sky130_fd_sc_hd__nand2_1
Xfanout79 _1147_ VGND VGND VDPWR VDPWR net79 sky130_fd_sc_hd__buf_2
Xfanout57 net59 VGND VGND VDPWR VDPWR net57 sky130_fd_sc_hd__buf_4
Xfanout68 net71 VGND VGND VDPWR VDPWR net68 sky130_fd_sc_hd__buf_2
Xfanout46 net47 VGND VGND VDPWR VDPWR net46 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_44_172 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_75_616 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[62\].gen_latches\[2\].p_latch net230 dig_ctrl_inst.latch_mem_inst.gclk\[62\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[62\]\[2\] sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_41_Left_119 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
Xclkload16 clknet_leaf_9_clk VGND VGND VDPWR VDPWR clkload16/Y sky130_fd_sc_hd__inv_12
Xdig_ctrl_inst.latch_mem_inst.gen_words\[51\].gen_latches\[0\].p_latch net241 dig_ctrl_inst.latch_mem_inst.gclk\[51\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[51\]\[0\] sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[19\].clock_buffer dig_ctrl_inst.latch_mem_inst.gen_gclk\[19\]._gclk
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.gclk\[19\] sky130_fd_sc_hd__clkbuf_4
X_1420_ net250 dig_ctrl_inst.spi_data_o\[5\] _1103_ _0162_ VGND VGND VDPWR VDPWR dig_ctrl_inst.data_out\[5\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_50_153 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_1351_ net151 _0132_ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.data_we\[31\]
+ sky130_fd_sc_hd__and2_1
X_1282_ _1076_ _1078_ net134 VGND VGND VDPWR VDPWR _1129_ sky130_fd_sc_hd__and3_4
XPHY_EDGE_ROW_50_Left_128 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
X_1618_ dig_ctrl_inst.latch_mem_inst.RAM\[17\]\[0\] _0120_ _0131_ dig_ctrl_inst.latch_mem_inst.RAM\[29\]\[0\]
+ VGND VGND VDPWR VDPWR _0330_ sky130_fd_sc_hd__a22o_1
XFILLER_0_26_183 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_81 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
Xfanout214 net323 VGND VGND VDPWR VDPWR net214 sky130_fd_sc_hd__buf_2
Xfanout247 net325 VGND VGND VDPWR VDPWR net247 sky130_fd_sc_hd__buf_1
Xfanout203 net207 VGND VGND VDPWR VDPWR net203 sky130_fd_sc_hd__clkbuf_2
Xfanout258 net259 VGND VGND VDPWR VDPWR net258 sky130_fd_sc_hd__buf_4
Xfanout236 net327 VGND VGND VDPWR VDPWR net236 sky130_fd_sc_hd__clkbuf_2
Xfanout225 net231 VGND VGND VDPWR VDPWR net225 sky130_fd_sc_hd__buf_2
X_1549_ _0245_ _0261_ _0253_ _0257_ VGND VGND VDPWR VDPWR _0262_ sky130_fd_sc_hd__or4b_1
XTAP_TAPCELL_ROW_37_384 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[48\].clock_gate clknet_leaf_12_clk dig_ctrl_inst.latch_mem_inst.data_we\[48\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.gen_gclk\[48\]._gclk sky130_fd_sc_hd__dlclkp_1
XTAP_TAPCELL_ROW_20_284 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_18 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_8
Xdig_ctrl_inst.latch_mem_inst.gen_words\[55\].gen_latches\[1\].p_latch net233 dig_ctrl_inst.latch_mem_inst.gclk\[55\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[55\]\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_55_256 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_223 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_309 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_6
X_2521_ net279 VGND VGND VDPWR VDPWR uio_oe[2] sky130_fd_sc_hd__buf_2
XFILLER_0_11_337 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_175 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_1403_ net153 _0156_ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.data_we\[59\]
+ sky130_fd_sc_hd__and2_1
X_2383_ clknet_leaf_4_clk net331 net174 VGND VGND VDPWR VDPWR dig_ctrl_inst.synchronizer_port_i_inst\[5\].out
+ sky130_fd_sc_hd__dfrtp_1
X_1334_ net95 net68 VGND VGND VDPWR VDPWR _0125_ sky130_fd_sc_hd__and2_1
X_1265_ net182 _1026_ _1027_ dig_ctrl_inst.cpu_inst.ip\[4\] VGND VGND VDPWR VDPWR
+ _1113_ sky130_fd_sc_hd__o211a_1
XPHY_EDGE_ROW_18_Right_18 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
X_2452_ clknet_leaf_11_clk _0060_ net140 VGND VGND VDPWR VDPWR dig_ctrl_inst.cpu_inst.r1\[7\]
+ sky130_fd_sc_hd__dfrtp_1
Xinput3 ui_in[0] VGND VGND VDPWR VDPWR net3 sky130_fd_sc_hd__clkbuf_1
X_1196_ net268 net264 dig_ctrl_inst.cpu_inst.r0\[3\] VGND VGND VDPWR VDPWR _1044_
+ sky130_fd_sc_hd__or3_1
XPHY_EDGE_ROW_27_Right_27 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[50\].clock_gate clknet_leaf_16_clk dig_ctrl_inst.latch_mem_inst.data_we\[50\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.gen_gclk\[50\]._gclk sky130_fd_sc_hd__dlclkp_1
XPHY_EDGE_ROW_36_Right_36 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[32\].gen_latches\[6\].p_latch net191 dig_ctrl_inst.latch_mem_inst.gclk\[32\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[32\]\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_69_337 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_45_Right_45 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_245 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[21\].gen_latches\[4\].p_latch net210 dig_ctrl_inst.latch_mem_inst.gclk\[21\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[21\]\[4\] sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_54_Right_54 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[59\].gen_latches\[2\].p_latch net230 dig_ctrl_inst.latch_mem_inst.gclk\[59\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[59\]\[2\] sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[10\].gen_latches\[2\].p_latch net228 dig_ctrl_inst.latch_mem_inst.gclk\[10\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[10\]\[2\] sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_63_Right_63 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
X_1952_ dig_ctrl_inst.latch_mem_inst.RAM\[23\]\[6\] net102 net100 net62 VGND VGND
+ VDPWR VDPWR _0658_ sky130_fd_sc_hd__and4_1
X_1883_ dig_ctrl_inst.latch_mem_inst.RAM\[46\]\[5\] net75 net55 VGND VGND VDPWR VDPWR
+ _0590_ sky130_fd_sc_hd__and3_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[48\].gen_latches\[0\].p_latch net241 dig_ctrl_inst.latch_mem_inst.gclk\[48\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[48\]\[0\] sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_72_Right_72 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
X_2504_ clknet_leaf_5_clk _0101_ net178 VGND VGND VDPWR VDPWR net34 sky130_fd_sc_hd__dfrtp_1
X_2435_ clknet_leaf_8_clk _0043_ VGND VGND VDPWR VDPWR dig_ctrl_inst.cpu_inst.prev_state\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_1248_ net251 dig_ctrl_inst.spi_receiver_inst.stb_o VGND VGND VDPWR VDPWR _1096_
+ sky130_fd_sc_hd__nand2_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[3\].gen_latches\[4\].p_latch net212 dig_ctrl_inst.latch_mem_inst.gclk\[3\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[3\]\[4\] sky130_fd_sc_hd__dlxtp_1
X_1317_ net123 net73 VGND VGND VDPWR VDPWR _0116_ sky130_fd_sc_hd__and2_1
X_2366_ _0685_ _0740_ _1009_ VGND VGND VDPWR VDPWR _0993_ sky130_fd_sc_hd__or3b_4
X_2297_ _0751_ _0964_ _0963_ VGND VGND VDPWR VDPWR _0975_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_2_41 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_329 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_82 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
X_1179_ net182 _1010_ VGND VGND VDPWR VDPWR _1027_ sky130_fd_sc_hd__or2_4
XANTENNA_30 dig_ctrl_inst.spi_data_i\[0\] VGND VGND VDPWR VDPWR sky130_fd_sc_hd__diode_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[36\].gen_latches\[7\].p_latch net185 dig_ctrl_inst.latch_mem_inst.gclk\[36\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[36\]\[7\] sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[25\].gen_latches\[5\].p_latch net203 dig_ctrl_inst.latch_mem_inst.gclk\[25\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[25\]\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_69_189 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
Xdig_ctrl_inst.latch_mem_inst.gen_input_latches\[5\].n_latch dig_ctrl_inst.data_out\[5\]
+ clknet_leaf_8_clk VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.wdata\[5\]
+ sky130_fd_sc_hd__dlxtn_1
XTAP_TAPCELL_ROW_53_482 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_204 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[14\].gen_latches\[3\].p_latch net220 dig_ctrl_inst.latch_mem_inst.gclk\[14\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[14\]\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_0_337 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
X_2082_ net160 net137 VGND VGND VDPWR VDPWR _0775_ sky130_fd_sc_hd__nand2_1
X_2220_ _1068_ _0776_ _0815_ VGND VGND VDPWR VDPWR _0908_ sky130_fd_sc_hd__o21ba_1
X_2151_ net166 net164 net161 VGND VGND VDPWR VDPWR _0842_ sky130_fd_sc_hd__or3_1
XFILLER_0_75_137 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_329 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
X_1866_ dig_ctrl_inst.latch_mem_inst.RAM\[38\]\[5\] net95 net59 VGND VGND VDPWR VDPWR
+ _0573_ sky130_fd_sc_hd__and3_2
X_1797_ dig_ctrl_inst.latch_mem_inst.RAM\[0\]\[3\] _0288_ net39 _0504_ VGND VGND VDPWR
+ VDPWR _0506_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_31_218 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_1935_ dig_ctrl_inst.latch_mem_inst.RAM\[57\]\[6\] net116 net90 net43 VGND VGND VDPWR
+ VDPWR _0641_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_59_519 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[7\].gen_latches\[5\].p_latch net206 dig_ctrl_inst.latch_mem_inst.gclk\[7\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[7\]\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_58_71 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
X_2418_ clknet_leaf_8_clk _0026_ net143 VGND VGND VDPWR VDPWR dig_ctrl_inst.cpu_inst.arg0\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_2349_ dig_ctrl_inst.cpu_inst.port_o\[4\] net32 _0987_ VGND VGND VDPWR VDPWR _0099_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_50_463 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_419 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_318 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_0_Right_0 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_262 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_29 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[29\].gen_latches\[6\].p_latch net197 dig_ctrl_inst.latch_mem_inst.gclk\[29\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[29\]\[6\] sky130_fd_sc_hd__dlxtp_1
Xhold108 net28 VGND VGND VDPWR VDPWR net390 sky130_fd_sc_hd__dlygate4sd3_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[18\].gen_latches\[4\].p_latch net213 dig_ctrl_inst.latch_mem_inst.gclk\[18\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[18\]\[4\] sky130_fd_sc_hd__dlxtp_1
X_1651_ dig_ctrl_inst.latch_mem_inst.RAM\[26\]\[1\] net294 net66 VGND VGND VDPWR VDPWR
+ _0362_ sky130_fd_sc_hd__and3_2
X_1720_ dig_ctrl_inst.latch_mem_inst.RAM\[23\]\[2\] _0126_ _0150_ dig_ctrl_inst.latch_mem_inst.RAM\[52\]\[2\]
+ VGND VGND VDPWR VDPWR _0430_ sky130_fd_sc_hd__a22o_1
X_1582_ dig_ctrl_inst.latch_mem_inst.RAM\[62\]\[0\] net73 net48 VGND VGND VDPWR VDPWR
+ _0294_ sky130_fd_sc_hd__and3_2
XFILLER_0_0_167 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_2065_ net300 _0755_ _0757_ _0199_ VGND VGND VDPWR VDPWR _0758_ sky130_fd_sc_hd__o211a_1
X_2203_ _0890_ _0891_ VGND VGND VDPWR VDPWR _0892_ sky130_fd_sc_hd__and2b_1
X_2134_ dig_ctrl_inst.cpu_inst.data\[1\] _0743_ _0825_ net164 VGND VGND VDPWR VDPWR
+ _0826_ sky130_fd_sc_hd__a22o_1
XFILLER_0_60_83 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_173 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_1849_ dig_ctrl_inst.latch_mem_inst.RAM\[1\]\[4\] _1130_ _0131_ dig_ctrl_inst.latch_mem_inst.RAM\[29\]\[4\]
+ VGND VGND VDPWR VDPWR _0557_ sky130_fd_sc_hd__a22o_1
X_1918_ dig_ctrl_inst.latch_mem_inst.RAM\[18\]\[6\] net111 net68 VGND VGND VDPWR VDPWR
+ _0624_ sky130_fd_sc_hd__and3_2
XFILLER_0_39_137 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_4_188 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_118 VDPWR VGND VDPWR VGND sky130_ef_sc_hd__decap_12
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[55\].clock_gate clknet_leaf_17_clk dig_ctrl_inst.latch_mem_inst.data_we\[55\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.gen_gclk\[55\]._gclk sky130_fd_sc_hd__dlclkp_1
XFILLER_0_53_162 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_140 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
X_1703_ dig_ctrl_inst.latch_mem_inst.RAM\[14\]\[2\] net123 net73 VGND VGND VDPWR VDPWR
+ _0413_ sky130_fd_sc_hd__and3_2
Xclkbuf_leaf_11_clk clknet_1_0__leaf_clk VGND VGND VDPWR VDPWR clknet_leaf_11_clk
+ sky130_fd_sc_hd__clkbuf_8
X_1634_ dig_ctrl_inst.latch_mem_inst.RAM\[61\]\[1\] net115 net80 net43 VGND VGND VDPWR
+ VDPWR _0345_ sky130_fd_sc_hd__and4_1
X_1565_ net125 net97 VGND VGND VDPWR VDPWR _0277_ sky130_fd_sc_hd__and2_2
X_1496_ _1060_ dig_ctrl_inst.cpu_inst.data\[2\] _0198_ VGND VGND VDPWR VDPWR _0213_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_76_221 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
X_2048_ dig_ctrl_inst.cpu_inst.cpu_state\[2\] net354 _0161_ VGND VGND VDPWR VDPWR
+ _0044_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_1_169 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2117_ _0258_ _0760_ _0766_ net157 VGND VGND VDPWR VDPWR _0809_ sky130_fd_sc_hd__o22a_1
XFILLER_0_12_3 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
Xfanout69 net71 VGND VGND VDPWR VDPWR net69 sky130_fd_sc_hd__buf_2
Xfanout58 net59 VGND VGND VDPWR VDPWR net58 sky130_fd_sc_hd__buf_2
Xfanout47 _0147_ VGND VGND VDPWR VDPWR net47 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_17_310 VDPWR VGND VDPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_617 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[62\].gen_latches\[6\].p_latch net195 dig_ctrl_inst.latch_mem_inst.gclk\[62\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[62\]\[6\] sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[58\].clock_buffer dig_ctrl_inst.latch_mem_inst.gen_gclk\[58\]._gclk
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.gclk\[58\] sky130_fd_sc_hd__clkbuf_4
Xclkload17 clknet_leaf_19_clk VGND VGND VDPWR VDPWR clkload17/Y sky130_fd_sc_hd__inv_12
Xdig_ctrl_inst.latch_mem_inst.gen_words\[51\].gen_latches\[4\].p_latch net212 dig_ctrl_inst.latch_mem_inst.gclk\[51\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[51\]\[4\] sky130_fd_sc_hd__dlxtp_1
X_1350_ net106 net82 net69 VGND VGND VDPWR VDPWR _0132_ sky130_fd_sc_hd__and3_4
X_1281_ net130 net152 net121 VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.data_we\[0\]
+ sky130_fd_sc_hd__and3_2
Xclkbuf_leaf_0_clk clknet_1_1__leaf_clk VGND VGND VDPWR VDPWR clknet_leaf_0_clk sky130_fd_sc_hd__clkbuf_8
Xdig_ctrl_inst.latch_mem_inst.gen_words\[40\].gen_latches\[2\].p_latch net224 dig_ctrl_inst.latch_mem_inst.gclk\[40\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[40\]\[2\] sky130_fd_sc_hd__dlxtp_1
Xfanout204 net206 VGND VGND VDPWR VDPWR net204 sky130_fd_sc_hd__clkbuf_2
X_1617_ dig_ctrl_inst.latch_mem_inst.RAM\[44\]\[0\] _0144_ _0148_ dig_ctrl_inst.latch_mem_inst.RAM\[49\]\[0\]
+ VGND VGND VDPWR VDPWR _0329_ sky130_fd_sc_hd__a22o_1
XFILLER_0_41_132 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_295 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_262 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
Xfanout237 net238 VGND VGND VDPWR VDPWR net237 sky130_fd_sc_hd__clkbuf_2
Xfanout248 dig_ctrl_inst.cpu_inst.cpu_state\[0\] VGND VGND VDPWR VDPWR net248 sky130_fd_sc_hd__clkbuf_4
Xfanout226 net227 VGND VGND VDPWR VDPWR net226 sky130_fd_sc_hd__clkbuf_2
Xfanout259 dig_ctrl_inst.cpu_inst.arg1\[0\] VGND VGND VDPWR VDPWR net259 sky130_fd_sc_hd__buf_2
Xfanout215 net216 VGND VGND VDPWR VDPWR net215 sky130_fd_sc_hd__clkbuf_2
X_1548_ _0258_ _0260_ VGND VGND VDPWR VDPWR _0261_ sky130_fd_sc_hd__and2_1
X_1479_ net285 _1031_ VGND VGND VDPWR VDPWR _0198_ sky130_fd_sc_hd__or2_2
XTAP_TAPCELL_ROW_37_385 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_154 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_285 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_3 VDPWR VGND VDPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_338 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_29 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_28_330 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[55\].gen_latches\[5\].p_latch net203 dig_ctrl_inst.latch_mem_inst.gclk\[55\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[55\]\[5\] sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_11_230 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2520_ net270 VGND VGND VDPWR VDPWR uio_oe[1] sky130_fd_sc_hd__buf_2
X_1402_ net107 net92 net49 VGND VGND VDPWR VDPWR _0156_ sky130_fd_sc_hd__and3_2
X_2451_ clknet_leaf_10_clk _0059_ net142 VGND VGND VDPWR VDPWR dig_ctrl_inst.cpu_inst.r1\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_11_55 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_165 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
Xinput4 ui_in[1] VGND VGND VDPWR VDPWR net4 sky130_fd_sc_hd__clkbuf_1
X_2382_ clknet_leaf_3_clk net8 net175 VGND VGND VDPWR VDPWR dig_ctrl_inst.synchronizer_port_i_inst\[5\].pipe\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[44\].gen_latches\[3\].p_latch net221 dig_ctrl_inst.latch_mem_inst.gclk\[44\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[44\]\[3\] sky130_fd_sc_hd__dlxtp_1
X_1264_ _1098_ _1105_ _1111_ dig_ctrl_inst.spi_addr\[5\] _1002_ VGND VGND VDPWR VDPWR
+ _1112_ sky130_fd_sc_hd__o32a_4
XFILLER_0_36_41 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_6
X_1333_ net150 _0124_ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.data_we\[21\]
+ sky130_fd_sc_hd__and2_1
X_1195_ net264 dig_ctrl_inst.cpu_inst.r1\[3\] VGND VGND VDPWR VDPWR _1043_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_34_366 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[33\].gen_latches\[1\].p_latch net233 dig_ctrl_inst.latch_mem_inst.gclk\[33\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[33\]\[1\] sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[10\].gen_latches\[6\].p_latch net195 dig_ctrl_inst.latch_mem_inst.gclk\[10\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[10\]\[6\] sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[59\].gen_latches\[6\].p_latch net195 dig_ctrl_inst.latch_mem_inst.gclk\[59\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[59\]\[6\] sky130_fd_sc_hd__dlxtp_1
X_1882_ dig_ctrl_inst.latch_mem_inst.RAM\[23\]\[5\] net103 net100 net63 VGND VGND
+ VDPWR VDPWR _0589_ sky130_fd_sc_hd__and4_1
X_1951_ dig_ctrl_inst.latch_mem_inst.RAM\[52\]\[6\] net96 net43 VGND VGND VDPWR VDPWR
+ _0657_ sky130_fd_sc_hd__and3_2
X_2503_ clknet_leaf_5_clk _0100_ net177 VGND VGND VDPWR VDPWR net33 sky130_fd_sc_hd__dfrtp_1
X_2434_ clknet_leaf_8_clk net347 VGND VGND VDPWR VDPWR dig_ctrl_inst.cpu_inst.prev_state\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_2365_ _0506_ _0565_ _0623_ VGND VGND VDPWR VDPWR _0992_ sky130_fd_sc_hd__and3_2
XFILLER_0_11_113 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[48\].gen_latches\[4\].p_latch net323 dig_ctrl_inst.latch_mem_inst.gclk\[48\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[48\]\[4\] sky130_fd_sc_hd__dlxtp_1
X_1316_ _1075_ _1077_ _1093_ net135 _1047_ VGND VGND VDPWR VDPWR _0115_ sky130_fd_sc_hd__o2111a_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[37\].gen_latches\[2\].p_latch net228 dig_ctrl_inst.latch_mem_inst.gclk\[37\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[37\]\[2\] sky130_fd_sc_hd__dlxtp_1
X_1247_ _1076_ _1078_ _1093_ net135 _1047_ VGND VGND VDPWR VDPWR _1095_ sky130_fd_sc_hd__a2111oi_1
X_2296_ net361 _0974_ _0967_ VGND VGND VDPWR VDPWR _0059_ sky130_fd_sc_hd__mux2_1
X_1178_ net298 _1019_ net283 _1015_ _1011_ VGND VGND VDPWR VDPWR _1026_ sky130_fd_sc_hd__o32ai_4
XFILLER_0_74_341 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XANTENNA_31 net19 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__diode_2
XANTENNA_20 net100 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__diode_2
XFILLER_0_2_97 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[26\].gen_latches\[0\].p_latch net246 dig_ctrl_inst.latch_mem_inst.gclk\[26\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[26\]\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_6_195 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_113 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_53_483 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[14\].gen_latches\[7\].p_latch net185 dig_ctrl_inst.latch_mem_inst.gclk\[14\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[14\]\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_0_305 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
X_2150_ _0838_ _0839_ _0840_ net167 net170 VGND VGND VDPWR VDPWR _0841_ sky130_fd_sc_hd__a221o_1
X_2081_ _0763_ _0765_ _0773_ VGND VGND VDPWR VDPWR _0774_ sky130_fd_sc_hd__o21a_1
XFILLER_0_17_54 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
X_1934_ dig_ctrl_inst.latch_mem_inst.RAM\[17\]\[6\] net132 net118 net68 VGND VGND
+ VDPWR VDPWR _0640_ sky130_fd_sc_hd__and4_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[8\].gen_latches\[0\].p_latch net242 dig_ctrl_inst.latch_mem_inst.gclk\[8\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[8\]\[0\] sky130_fd_sc_hd__dlxtp_1
X_1865_ dig_ctrl_inst.latch_mem_inst.RAM\[10\]\[5\] net124 net83 VGND VGND VDPWR VDPWR
+ _0572_ sky130_fd_sc_hd__and3_2
X_1796_ net39 _0504_ dig_ctrl_inst.latch_mem_inst.RAM\[0\]\[3\] _0288_ VGND VGND VDPWR
+ VDPWR _0505_ sky130_fd_sc_hd__o2bb2a_1
X_2348_ dig_ctrl_inst.cpu_inst.port_o\[3\] net31 _0987_ VGND VGND VDPWR VDPWR _0098_
+ sky130_fd_sc_hd__mux2_1
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[62\].clock_gate clknet_leaf_0_clk dig_ctrl_inst.latch_mem_inst.data_we\[62\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.gen_gclk\[62\]._gclk sky130_fd_sc_hd__dlclkp_1
XFILLER_0_42_3 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_2417_ clknet_leaf_10_clk _0025_ net140 VGND VGND VDPWR VDPWR dig_ctrl_inst.cpu_inst.skip
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_10_Left_88 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_67_564 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2279_ dig_ctrl_inst.synchronizer_port_i_inst\[7\].out _0802_ _0804_ dig_ctrl_inst.spi_data_o\[7\]
+ VGND VGND VDPWR VDPWR _0965_ sky130_fd_sc_hd__a22oi_2
XTAP_TAPCELL_ROW_50_464 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_341 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_219 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_341 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
Xhold109 dig_ctrl_inst.spi_receiver_inst.spi_cnt\[2\] VGND VGND VDPWR VDPWR net391
+ sky130_fd_sc_hd__dlygate4sd3_1
X_1581_ dig_ctrl_inst.latch_mem_inst.RAM\[61\]\[0\] net118 net82 net48 VGND VGND VDPWR
+ VDPWR _0293_ sky130_fd_sc_hd__and4_1
XFILLER_0_53_333 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
X_1650_ dig_ctrl_inst.latch_mem_inst.RAM\[50\]\[1\] net109 net42 VGND VGND VDPWR VDPWR
+ _0361_ sky130_fd_sc_hd__and3_2
X_2202_ net159 _0867_ VGND VGND VDPWR VDPWR _0891_ sky130_fd_sc_hd__nand2_1
XFILLER_0_0_113 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_146 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_85 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_41 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
X_2064_ _1020_ _1024_ _0756_ VGND VGND VDPWR VDPWR _0757_ sky130_fd_sc_hd__a21o_1
X_2133_ _1015_ _1019_ VGND VGND VDPWR VDPWR _0825_ sky130_fd_sc_hd__nor2_2
XFILLER_0_29_341 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_1917_ net252 _0622_ _0276_ VGND VGND VDPWR VDPWR _0031_ sky130_fd_sc_hd__mux2_1
XFILLER_0_69_93 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_71 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[8\].clock_buffer dig_ctrl_inst.latch_mem_inst.gen_gclk\[8\]._gclk
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.gclk\[8\] sky130_fd_sc_hd__clkbuf_4
X_1848_ dig_ctrl_inst.latch_mem_inst.RAM\[9\]\[4\] _1143_ _0155_ dig_ctrl_inst.latch_mem_inst.RAM\[58\]\[4\]
+ VGND VGND VDPWR VDPWR _0556_ sky130_fd_sc_hd__a22o_1
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[22\].clock_buffer dig_ctrl_inst.latch_mem_inst.gen_gclk\[22\]._gclk
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.gclk\[22\] sky130_fd_sc_hd__clkbuf_4
X_1779_ dig_ctrl_inst.latch_mem_inst.RAM\[46\]\[3\] net72 net56 VGND VGND VDPWR VDPWR
+ _0488_ sky130_fd_sc_hd__and3_2
XTAP_TAPCELL_ROW_4_189 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_141 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_160 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
X_1564_ net182 _0200_ VGND VGND VDPWR VDPWR _0276_ sky130_fd_sc_hd__and2_2
X_1633_ dig_ctrl_inst.latch_mem_inst.RAM\[59\]\[1\] net102 net90 net42 VGND VGND VDPWR
+ VDPWR _0344_ sky130_fd_sc_hd__and4_1
X_1702_ dig_ctrl_inst.latch_mem_inst.RAM\[48\]\[2\] net130 net46 VGND VGND VDPWR VDPWR
+ _0412_ sky130_fd_sc_hd__and3_2
X_1495_ dig_ctrl_inst.cpu_inst.ip\[0\] dig_ctrl_inst.cpu_inst.ip\[1\] _0210_ VGND
+ VGND VDPWR VDPWR _0212_ sky130_fd_sc_hd__and3_2
X_2047_ dig_ctrl_inst.cpu_inst.cpu_state\[1\] net349 _0161_ VGND VGND VDPWR VDPWR
+ _0043_ sky130_fd_sc_hd__mux2_1
X_2116_ _0761_ _0776_ net157 VGND VGND VDPWR VDPWR _0808_ sky130_fd_sc_hd__mux2_1
Xfanout48 net49 VGND VGND VDPWR VDPWR net48 sky130_fd_sc_hd__buf_4
Xfanout59 net60 VGND VGND VDPWR VDPWR net59 sky130_fd_sc_hd__buf_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[63\].gen_latches\[1\].p_latch net237 dig_ctrl_inst.latch_mem_inst.gclk\[63\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[63\]\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_44_141 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_322 VDPWR VGND VDPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_282 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_13_Left_91 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_108 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
X_1280_ _1112_ _1127_ VGND VGND VDPWR VDPWR _1128_ sky130_fd_sc_hd__nor2_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[40\].gen_latches\[6\].p_latch net196 dig_ctrl_inst.latch_mem_inst.gclk\[40\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[40\]\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_25_10 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_43 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_54 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_75 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_42 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_14_250 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout205 net206 VGND VGND VDPWR VDPWR net205 sky130_fd_sc_hd__buf_1
X_1616_ dig_ctrl_inst.latch_mem_inst.RAM\[19\]\[0\] _0122_ _0293_ _0294_ _0302_ VGND
+ VGND VDPWR VDPWR _0328_ sky130_fd_sc_hd__a2111o_1
Xfanout238 net239 VGND VGND VDPWR VDPWR net238 sky130_fd_sc_hd__clkbuf_2
Xfanout227 net231 VGND VGND VDPWR VDPWR net227 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_5_31 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_8
X_1547_ net158 net164 VGND VGND VDPWR VDPWR _0260_ sky130_fd_sc_hd__or2_1
Xfanout216 net329 VGND VGND VDPWR VDPWR net216 sky130_fd_sc_hd__buf_2
X_1478_ dig_ctrl_inst.cpu_inst.r0\[7\] dig_ctrl_inst.cpu_inst.port_o\[7\] _0176_ VGND
+ VGND VDPWR VDPWR _0018_ sky130_fd_sc_hd__mux2_1
Xfanout249 net251 VGND VGND VDPWR VDPWR net249 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_49_222 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_37_386 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_341 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_286 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_317 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[56\].gen_latches\[0\].p_latch net242 dig_ctrl_inst.latch_mem_inst.gclk\[56\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[56\]\[0\] sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_28_331 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_231 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1401_ net155 net85 net50 VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.data_we\[58\]
+ sky130_fd_sc_hd__and3_2
X_2381_ clknet_leaf_4_clk net338 net174 VGND VGND VDPWR VDPWR dig_ctrl_inst.synchronizer_port_i_inst\[6\].out
+ sky130_fd_sc_hd__dfrtp_1
X_2450_ clknet_leaf_7_clk _0058_ net144 VGND VGND VDPWR VDPWR dig_ctrl_inst.cpu_inst.r1\[5\]
+ sky130_fd_sc_hd__dfrtp_1
Xinput5 ui_in[2] VGND VGND VDPWR VDPWR net5 sky130_fd_sc_hd__clkbuf_1
X_1194_ net267 dig_ctrl_inst.cpu_inst.r2\[3\] VGND VGND VDPWR VDPWR _1042_ sky130_fd_sc_hd__and2b_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[44\].gen_latches\[7\].p_latch net189 dig_ctrl_inst.latch_mem_inst.gclk\[44\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[44\]\[7\] sky130_fd_sc_hd__dlxtp_1
X_1263_ _1039_ _1110_ net249 VGND VGND VDPWR VDPWR _1111_ sky130_fd_sc_hd__a21o_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[0\].gen_latches\[2\].p_latch net226 dig_ctrl_inst.latch_mem_inst.gclk\[0\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[0\]\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_36_75 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_1332_ net116 net99 net62 VGND VGND VDPWR VDPWR _0124_ sky130_fd_sc_hd__and3_2
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[15\].clock_buffer dig_ctrl_inst.latch_mem_inst.gen_gclk\[15\]._gclk
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.gclk\[15\] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_52_85 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_34_367 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_3 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_291 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_280 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[33\].gen_latches\[5\].p_latch net201 dig_ctrl_inst.latch_mem_inst.gclk\[33\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[33\]\[5\] sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[22\].gen_latches\[3\].p_latch net220 dig_ctrl_inst.latch_mem_inst.gclk\[22\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[22\]\[3\] sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_25_312 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[11\].gen_latches\[1\].p_latch net238 dig_ctrl_inst.latch_mem_inst.gclk\[11\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[11\]\[1\] sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_29_Left_107 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
X_1950_ dig_ctrl_inst.latch_mem_inst.RAM\[40\]\[6\] net88 net57 VGND VGND VDPWR VDPWR
+ _0656_ sky130_fd_sc_hd__and3_2
XPHY_EDGE_ROW_38_Left_116 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_22 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_6
X_2502_ clknet_leaf_5_clk _0099_ net177 VGND VGND VDPWR VDPWR net32 sky130_fd_sc_hd__dfrtp_1
X_1881_ dig_ctrl_inst.latch_mem_inst.RAM\[1\]\[5\] _1130_ _0152_ dig_ctrl_inst.latch_mem_inst.RAM\[54\]\[5\]
+ _0587_ VGND VGND VDPWR VDPWR _0588_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_31_348 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_325 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_77 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_99 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
X_1315_ net155 _0114_ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.data_we\[13\]
+ sky130_fd_sc_hd__and2_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[4\].gen_latches\[3\].p_latch net220 dig_ctrl_inst.latch_mem_inst.gclk\[4\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[4\]\[3\] sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_47_Left_125 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
X_2364_ _0338_ _0398_ _0506_ _0623_ VGND VGND VDPWR VDPWR _0991_ sky130_fd_sc_hd__o211ai_1
X_2433_ clknet_leaf_13_clk _0041_ net139 VGND VGND VDPWR VDPWR dig_ctrl_inst.cpu_inst.data\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_56_Left_134 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
X_1246_ net249 _1079_ _1091_ _1085_ _1092_ VGND VGND VDPWR VDPWR _1094_ sky130_fd_sc_hd__o41ai_2
X_2295_ _0751_ _0946_ _0943_ VGND VGND VDPWR VDPWR _0974_ sky130_fd_sc_hd__o21ai_1
X_1177_ net181 _1019_ _1017_ _1015_ _1011_ VGND VGND VDPWR VDPWR _1025_ sky130_fd_sc_hd__o32a_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[37\].gen_latches\[6\].p_latch net195 dig_ctrl_inst.latch_mem_inst.gclk\[37\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[37\]\[6\] sky130_fd_sc_hd__dlxtp_1
XANTENNA_32 _1135_ VGND VGND VDPWR VDPWR sky130_fd_sc_hd__diode_2
XANTENNA_21 net329 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__diode_2
XANTENNA_10 dig_ctrl_inst.latch_mem_inst.gclk\[19\] VGND VGND VDPWR VDPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_65_Left_143 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_291 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_74_Left_152 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[26\].gen_latches\[4\].p_latch net211 dig_ctrl_inst.latch_mem_inst.gclk\[26\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[26\]\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_69_169 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_147 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
Xmax_cap89 _1141_ VGND VGND VDPWR VDPWR net89 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_53_484 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[15\].gen_latches\[2\].p_latch net229 dig_ctrl_inst.latch_mem_inst.gclk\[15\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[15\]\[2\] sky130_fd_sc_hd__dlxtp_1
X_2080_ _0767_ _0768_ _0771_ _0772_ VGND VGND VDPWR VDPWR _0773_ sky130_fd_sc_hd__o211a_1
XFILLER_0_17_11 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_65 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_1933_ dig_ctrl_inst.latch_mem_inst.RAM\[12\]\[6\] net122 net76 VGND VGND VDPWR VDPWR
+ _0639_ sky130_fd_sc_hd__and3_2
X_1864_ dig_ctrl_inst.latch_mem_inst.RAM\[56\]\[5\] net88 net49 VGND VGND VDPWR VDPWR
+ _0571_ sky130_fd_sc_hd__and3_2
X_1795_ _0464_ _0469_ _0486_ _0503_ VGND VGND VDPWR VDPWR _0504_ sky130_fd_sc_hd__nor4_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[8\].gen_latches\[4\].p_latch net209 dig_ctrl_inst.latch_mem_inst.gclk\[8\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[8\]\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_24_250 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
X_2347_ dig_ctrl_inst.cpu_inst.port_o\[2\] net30 _0987_ VGND VGND VDPWR VDPWR _0097_
+ sky130_fd_sc_hd__mux2_1
X_2278_ _0233_ _0944_ VGND VGND VDPWR VDPWR _0964_ sky130_fd_sc_hd__xor2_1
X_2416_ clknet_leaf_13_clk _0024_ net140 VGND VGND VDPWR VDPWR dig_ctrl_inst.cpu_inst.ip\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_66_139 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_67_565 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1229_ dig_ctrl_inst.spi_addr\[0\] _1002_ VGND VGND VDPWR VDPWR _1077_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_50_465 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_510 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[19\].gen_latches\[3\].p_latch net215 dig_ctrl_inst.latch_mem_inst.gclk\[19\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[19\]\[3\] sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_41_410 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1580_ dig_ctrl_inst.latch_mem_inst.RAM\[24\]\[0\] net87 net66 VGND VGND VDPWR VDPWR
+ _0292_ sky130_fd_sc_hd__and3_2
XFILLER_0_0_103 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_8
X_2201_ net159 _0867_ VGND VGND VDPWR VDPWR _0890_ sky130_fd_sc_hd__nor2_1
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[61\].clock_buffer dig_ctrl_inst.latch_mem_inst.gen_gclk\[61\]._gclk
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.gclk\[61\] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_0_169 VDPWR VGND VDPWR VGND sky130_ef_sc_hd__decap_12
X_2132_ _0255_ _0785_ _0793_ _0254_ _0823_ VGND VGND VDPWR VDPWR _0824_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_64_546 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_139 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_2063_ _0751_ _0753_ VGND VGND VDPWR VDPWR _0756_ sky130_fd_sc_hd__or2_4
X_1847_ dig_ctrl_inst.latch_mem_inst.RAM\[59\]\[4\] _0156_ _0552_ _0553_ _0554_ VGND
+ VGND VDPWR VDPWR _0555_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_63_109 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
X_1916_ dig_ctrl_inst.latch_mem_inst.RAM\[0\]\[5\] _0288_ net37 net36 VGND VGND VDPWR
+ VDPWR _0623_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_71_186 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_253 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
X_1778_ dig_ctrl_inst.latch_mem_inst.RAM\[32\]\[3\] net129 net56 VGND VGND VDPWR VDPWR
+ _0487_ sky130_fd_sc_hd__and3_2
XFILLER_0_35_312 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
X_1701_ dig_ctrl_inst.latch_mem_inst.RAM\[50\]\[2\] net111 net50 VGND VGND VDPWR VDPWR
+ _0411_ sky130_fd_sc_hd__and3_2
X_2523__272 VGND VGND VDPWR VDPWR _2523__272/HI net272 sky130_fd_sc_hd__conb_1
XFILLER_0_41_337 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_20 VDPWR VGND VDPWR VGND sky130_ef_sc_hd__decap_12
X_1494_ _0204_ _0210_ VGND VGND VDPWR VDPWR _0211_ sky130_fd_sc_hd__or2_1
X_1632_ dig_ctrl_inst.latch_mem_inst.RAM\[22\]\[1\] net94 net67 VGND VGND VDPWR VDPWR
+ _0343_ sky130_fd_sc_hd__and3_2
X_1563_ dig_ctrl_inst.cpu_inst.skip _0174_ _0274_ _0275_ VGND VGND VDPWR VDPWR _0025_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_55_63 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_2115_ dig_ctrl_inst.cpu_inst.r0\[0\] _0807_ net41 VGND VGND VDPWR VDPWR _0045_ sky130_fd_sc_hd__mux2_1
X_2530__276 VGND VGND VDPWR VDPWR _2530__276/HI net276 sky130_fd_sc_hd__conb_1
Xfanout49 net50 VGND VGND VDPWR VDPWR net49 sky130_fd_sc_hd__buf_4
X_2046_ dig_ctrl_inst.cpu_inst.cpu_state\[0\] net346 _0161_ VGND VGND VDPWR VDPWR
+ _0042_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_109 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_301 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_197 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_9_216 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_334 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[63\].gen_latches\[5\].p_latch net203 dig_ctrl_inst.latch_mem_inst.gclk\[63\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[63\]\[5\] sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_0_160 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_120 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[52\].gen_latches\[3\].p_latch net216 dig_ctrl_inst.latch_mem_inst.gclk\[52\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[52\]\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_76_29 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_175 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_337 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[41\].gen_latches\[1\].p_latch net236 dig_ctrl_inst.latch_mem_inst.gclk\[41\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[41\]\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_41_167 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_197 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_153 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_14_251 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1477_ dig_ctrl_inst.cpu_inst.r0\[6\] dig_ctrl_inst.cpu_inst.port_o\[6\] _0176_ VGND
+ VGND VDPWR VDPWR _0017_ sky130_fd_sc_hd__mux2_1
Xfanout239 net327 VGND VGND VDPWR VDPWR net239 sky130_fd_sc_hd__clkbuf_2
Xfanout206 net207 VGND VGND VDPWR VDPWR net206 sky130_fd_sc_hd__buf_1
Xfanout228 net231 VGND VGND VDPWR VDPWR net228 sky130_fd_sc_hd__clkbuf_2
X_1615_ dig_ctrl_inst.latch_mem_inst.RAM\[12\]\[0\] _1148_ _0278_ dig_ctrl_inst.latch_mem_inst.RAM\[5\]\[0\]
+ _0289_ VGND VGND VDPWR VDPWR _0327_ sky130_fd_sc_hd__a221o_1
XFILLER_0_41_189 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
Xfanout217 net219 VGND VGND VDPWR VDPWR net217 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_1_275 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
X_1546_ net158 net164 VGND VGND VDPWR VDPWR _0259_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_37_387 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2029_ _0730_ _0731_ _0732_ _0733_ VGND VGND VDPWR VDPWR _0734_ sky130_fd_sc_hd__or4_4
XTAP_TAPCELL_ROW_20_287 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[56\].gen_latches\[4\].p_latch net214 dig_ctrl_inst.latch_mem_inst.gclk\[56\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[56\]\[4\] sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_28_332 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_46 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_57 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_11_232 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[45\].gen_latches\[2\].p_latch net224 dig_ctrl_inst.latch_mem_inst.gclk\[45\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[45\]\[2\] sky130_fd_sc_hd__dlxtp_1
X_2380_ clknet_leaf_3_clk net9 net175 VGND VGND VDPWR VDPWR dig_ctrl_inst.synchronizer_port_i_inst\[6\].pipe\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_1400_ net83 _0147_ VGND VGND VDPWR VDPWR _0155_ sky130_fd_sc_hd__and2_2
X_1331_ net156 net97 net68 VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.data_we\[20\]
+ sky130_fd_sc_hd__and3_2
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[54\].clock_buffer dig_ctrl_inst.latch_mem_inst.gen_gclk\[54\]._gclk
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.gclk\[54\] sky130_fd_sc_hd__clkbuf_4
Xinput6 ui_in[3] VGND VGND VDPWR VDPWR net6 sky130_fd_sc_hd__clkbuf_1
X_1193_ net267 net264 dig_ctrl_inst.cpu_inst.r3\[3\] VGND VGND VDPWR VDPWR _1041_
+ sky130_fd_sc_hd__and3_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[34\].gen_latches\[0\].p_latch net245 dig_ctrl_inst.latch_mem_inst.gclk\[34\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[34\]\[0\] sky130_fd_sc_hd__dlxtp_1
X_1262_ net181 _1106_ _1107_ _1108_ _1109_ VGND VGND VDPWR VDPWR _1110_ sky130_fd_sc_hd__o41a_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[0\].gen_latches\[6\].p_latch net193 dig_ctrl_inst.latch_mem_inst.gclk\[0\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[0\]\[6\] sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_34_368 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_323 VDPWR VGND VDPWR VGND sky130_ef_sc_hd__decap_12
X_1529_ _1103_ net160 VGND VGND VDPWR VDPWR _0242_ sky130_fd_sc_hd__nand2_1
XFILLER_0_77_340 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[22\].gen_latches\[7\].p_latch net184 dig_ctrl_inst.latch_mem_inst.gclk\[22\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[22\]\[7\] sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_25_313 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_281 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_14_Right_14 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[11\].gen_latches\[5\].p_latch net204 dig_ctrl_inst.latch_mem_inst.gclk\[11\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[11\]\[5\] sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_23_Right_23 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_32_Right_32 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_31_349 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1880_ dig_ctrl_inst.latch_mem_inst.RAM\[40\]\[5\] net86 net60 VGND VGND VDPWR VDPWR
+ _0587_ sky130_fd_sc_hd__and3_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[49\].gen_latches\[3\].p_latch net217 dig_ctrl_inst.latch_mem_inst.gclk\[49\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[49\]\[3\] sky130_fd_sc_hd__dlxtp_1
X_2501_ clknet_leaf_5_clk _0098_ net178 VGND VGND VDPWR VDPWR net31 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_337 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[4\].gen_latches\[7\].p_latch net187 dig_ctrl_inst.latch_mem_inst.gclk\[4\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[4\]\[7\] sky130_fd_sc_hd__dlxtp_1
X_1314_ net126 net119 net82 VGND VGND VDPWR VDPWR _0114_ sky130_fd_sc_hd__and3_4
X_2294_ net365 _0973_ _0967_ VGND VGND VDPWR VDPWR _0058_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_41_Right_41 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
X_2363_ _0201_ _0989_ VGND VGND VDPWR VDPWR _0990_ sky130_fd_sc_hd__nand2_1
X_2432_ clknet_leaf_13_clk _0040_ net139 VGND VGND VDPWR VDPWR dig_ctrl_inst.cpu_inst.data\[6\]
+ sky130_fd_sc_hd__dfrtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[38\].gen_latches\[1\].p_latch net234 dig_ctrl_inst.latch_mem_inst.gclk\[38\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[38\]\[1\] sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_50_Right_50 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
X_1245_ net249 net289 _1091_ _1085_ _1092_ VGND VGND VDPWR VDPWR _1093_ sky130_fd_sc_hd__o41a_4
X_1176_ _0998_ net264 VGND VGND VDPWR VDPWR _1024_ sky130_fd_sc_hd__and2_1
XANTENNA_33 dig_ctrl_inst.cpu_inst.port_o\[5\] VGND VGND VDPWR VDPWR sky130_fd_sc_hd__diode_2
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[13\].clock_gate clknet_leaf_2_clk dig_ctrl_inst.latch_mem_inst.data_we\[13\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.gen_gclk\[13\]._gclk sky130_fd_sc_hd__dlclkp_1
XANTENNA_11 dig_ctrl_inst.latch_mem_inst.gclk\[32\] VGND VGND VDPWR VDPWR sky130_fd_sc_hd__diode_2
XANTENNA_22 net322 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__diode_2
XFILLER_0_42_251 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_192 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_53_485 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[15\].gen_latches\[6\].p_latch net191 dig_ctrl_inst.latch_mem_inst.gclk\[15\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[15\]\[6\] sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_44_430 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1932_ dig_ctrl_inst.latch_mem_inst.RAM\[10\]\[6\] net124 net83 VGND VGND VDPWR VDPWR
+ _0638_ sky130_fd_sc_hd__and3_2
X_1863_ dig_ctrl_inst.latch_mem_inst.RAM\[27\]\[5\] _0130_ _0278_ dig_ctrl_inst.latch_mem_inst.RAM\[5\]\[5\]
+ _0569_ VGND VGND VDPWR VDPWR _0570_ sky130_fd_sc_hd__a221o_1
XFILLER_0_33_99 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_2526__281 VGND VGND VDPWR VDPWR net281 _2526__281/LO sky130_fd_sc_hd__conb_1
X_1794_ _0490_ _0494_ _0498_ _0502_ VGND VGND VDPWR VDPWR _0503_ sky130_fd_sc_hd__or4_1
X_2415_ clknet_leaf_13_clk _0023_ net140 VGND VGND VDPWR VDPWR dig_ctrl_inst.cpu_inst.ip\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_2346_ dig_ctrl_inst.cpu_inst.port_o\[1\] net389 _0987_ VGND VGND VDPWR VDPWR _0096_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_67_566 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_85 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
X_1228_ dig_ctrl_inst.cpu_inst.ip\[0\] _1028_ _1067_ _1030_ _1074_ VGND VGND VDPWR
+ VDPWR _1076_ sky130_fd_sc_hd__a221o_2
XFILLER_0_28_3 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
X_2277_ _0788_ _0951_ _0962_ VGND VGND VDPWR VDPWR _0963_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_50_466 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_511 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[19\].gen_latches\[7\].p_latch net188 dig_ctrl_inst.latch_mem_inst.gclk\[19\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[19\]\[7\] sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_41_411 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[47\].clock_buffer dig_ctrl_inst.latch_mem_inst.gen_gclk\[47\]._gclk
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.gclk\[47\] sky130_fd_sc_hd__clkbuf_4
X_2062_ _0751_ _0753_ VGND VGND VDPWR VDPWR _0755_ sky130_fd_sc_hd__nor2_1
X_2200_ net167 _0771_ _0781_ _0888_ net170 VGND VGND VDPWR VDPWR _0889_ sky130_fd_sc_hd__a221o_1
X_2131_ _0786_ _0791_ net163 VGND VGND VDPWR VDPWR _0823_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_64_547 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_98 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_9 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_1846_ dig_ctrl_inst.latch_mem_inst.RAM\[56\]\[4\] net88 net49 VGND VGND VDPWR VDPWR
+ _0554_ sky130_fd_sc_hd__and3_2
XFILLER_0_60_97 VDPWR VGND VDPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_195 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_1915_ net37 net36 dig_ctrl_inst.latch_mem_inst.RAM\[0\]\[5\] _0288_ VGND VGND VDPWR
+ VDPWR _0622_ sky130_fd_sc_hd__o2bb2a_1
X_1777_ _0473_ _0477_ _0481_ _0485_ VGND VGND VDPWR VDPWR _0486_ sky130_fd_sc_hd__or4_1
XPHY_EDGE_ROW_4_Right_4 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
X_2329_ dig_ctrl_inst.spi_data_o\[1\] dig_ctrl_inst.spi_data_o\[2\] _0180_ VGND VGND
+ VDPWR VDPWR _0081_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_132 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_184 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_129 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
Xclone12 _1144_ VGND VGND VDPWR VDPWR net294 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_61_528 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_180 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1700_ dig_ctrl_inst.latch_mem_inst.RAM\[58\]\[2\] net85 net49 VGND VGND VDPWR VDPWR
+ _0410_ sky130_fd_sc_hd__and3_2
XFILLER_0_53_110 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_89 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_34 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_23 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_218 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_1631_ dig_ctrl_inst.latch_mem_inst.RAM\[28\]\[1\] net76 net67 VGND VGND VDPWR VDPWR
+ _0342_ sky130_fd_sc_hd__and3_2
Xclkbuf_leaf_3_clk clknet_1_1__leaf_clk VGND VGND VDPWR VDPWR clknet_leaf_3_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_39_32 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_6
X_1493_ dig_ctrl_inst.cpu_inst.ip\[0\] dig_ctrl_inst.cpu_inst.ip\[1\] dig_ctrl_inst.cpu_inst.ip\[2\]
+ _0173_ VGND VGND VDPWR VDPWR _0210_ sky130_fd_sc_hd__a31oi_1
X_1562_ dig_ctrl_inst.cpu_inst.instr\[6\] dig_ctrl_inst.cpu_inst.instr\[7\] _0175_
+ VGND VGND VDPWR VDPWR _0275_ sky130_fd_sc_hd__and3_2
XFILLER_0_55_53 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
X_2114_ _0798_ _0806_ VGND VGND VDPWR VDPWR _0807_ sky130_fd_sc_hd__nand2_1
X_2045_ net387 _0740_ _0741_ VGND VGND VDPWR VDPWR _0041_ sky130_fd_sc_hd__mux2_1
X_1829_ dig_ctrl_inst.latch_mem_inst.RAM\[41\]\[4\] net114 net90 net51 VGND VGND VDPWR
+ VDPWR _0537_ sky130_fd_sc_hd__and4_1
XFILLER_0_4_251 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_217 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[4\].clock_buffer dig_ctrl_inst.latch_mem_inst.gen_gclk\[4\]._gclk
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.gclk\[4\] sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_0_161 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_110 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[52\].gen_latches\[7\].p_latch net190 dig_ctrl_inst.latch_mem_inst.gclk\[52\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[52\]\[7\] sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[41\].gen_latches\[5\].p_latch net199 dig_ctrl_inst.latch_mem_inst.gclk\[41\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[41\]\[5\] sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[30\].gen_latches\[3\].p_latch net222 dig_ctrl_inst.latch_mem_inst.gclk\[30\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[30\]\[3\] sky130_fd_sc_hd__dlxtp_1
X_1614_ _0313_ _0318_ _0325_ VGND VGND VDPWR VDPWR _0326_ sky130_fd_sc_hd__or3_1
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[18\].clock_gate clknet_leaf_17_clk dig_ctrl_inst.latch_mem_inst.data_we\[18\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.gen_gclk\[18\]._gclk sky130_fd_sc_hd__dlclkp_1
XFILLER_0_66_85 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
Xfanout229 net230 VGND VGND VDPWR VDPWR net229 sky130_fd_sc_hd__clkbuf_2
X_1476_ dig_ctrl_inst.cpu_inst.r0\[5\] dig_ctrl_inst.cpu_inst.port_o\[5\] _0176_ VGND
+ VGND VDPWR VDPWR _0016_ sky130_fd_sc_hd__mux2_1
Xfanout207 net326 VGND VGND VDPWR VDPWR net207 sky130_fd_sc_hd__clkbuf_2
Xfanout218 net219 VGND VGND VDPWR VDPWR net218 sky130_fd_sc_hd__buf_1
X_1545_ dig_ctrl_inst.cpu_inst.r0\[0\] _1019_ _1065_ _1066_ net165 VGND VGND VDPWR
+ VDPWR _0258_ sky130_fd_sc_hd__o221ai_4
XFILLER_0_5_99 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_55 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_11 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_254 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_37_388 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_3 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
X_2028_ dig_ctrl_inst.latch_mem_inst.RAM\[13\]\[7\] _0114_ _0149_ dig_ctrl_inst.latch_mem_inst.RAM\[51\]\[7\]
+ VGND VGND VDPWR VDPWR _0733_ sky130_fd_sc_hd__a22o_1
XFILLER_0_17_165 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[20\].clock_gate clknet_leaf_19_clk dig_ctrl_inst.latch_mem_inst.data_we\[20\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.gen_gclk\[20\]._gclk sky130_fd_sc_hd__dlclkp_1
XTAP_TAPCELL_ROW_28_333 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_233 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[1\].gen_latches\[1\].p_latch net237 dig_ctrl_inst.latch_mem_inst.gclk\[1\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[1\]\[1\] sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[45\].gen_latches\[6\].p_latch net197 dig_ctrl_inst.latch_mem_inst.gclk\[45\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[45\]\[6\] sky130_fd_sc_hd__dlxtp_1
X_1330_ net97 net68 VGND VGND VDPWR VDPWR _0123_ sky130_fd_sc_hd__and2_1
X_1261_ net267 net263 dig_ctrl_inst.cpu_inst.r0\[5\] VGND VGND VDPWR VDPWR _1109_
+ sky130_fd_sc_hd__or3_1
Xinput7 ui_in[4] VGND VGND VDPWR VDPWR net7 sky130_fd_sc_hd__clkbuf_1
X_1192_ net248 dig_ctrl_inst.cpu_inst.cpu_state\[1\] _0999_ VGND VGND VDPWR VDPWR
+ _1040_ sky130_fd_sc_hd__or3_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[34\].gen_latches\[4\].p_latch net213 dig_ctrl_inst.latch_mem_inst.gclk\[34\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[34\]\[4\] sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_34_369 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_313 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_335 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_341 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[23\].gen_latches\[2\].p_latch net225 dig_ctrl_inst.latch_mem_inst.gclk\[23\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[23\]\[2\] sky130_fd_sc_hd__dlxtp_1
X_1459_ dig_ctrl_inst.spi_addr\[0\] dig_ctrl_inst.spi_addr\[1\] _0185_ dig_ctrl_inst.spi_addr\[2\]
+ VGND VGND VDPWR VDPWR _0190_ sky130_fd_sc_hd__a31o_1
X_1528_ _1103_ net160 VGND VGND VDPWR VDPWR _0241_ sky130_fd_sc_hd__and2_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[12\].gen_latches\[0\].p_latch net243 dig_ctrl_inst.latch_mem_inst.gclk\[12\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[12\]\[0\] sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_25_314 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_173 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[49\].gen_latches\[7\].p_latch net189 dig_ctrl_inst.latch_mem_inst.gclk\[49\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[49\]\[7\] sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[5\].gen_latches\[2\].p_latch net228 dig_ctrl_inst.latch_mem_inst.gclk\[5\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[5\]\[2\] sky130_fd_sc_hd__dlxtp_1
X_2500_ clknet_leaf_5_clk _0097_ net177 VGND VGND VDPWR VDPWR net30 sky130_fd_sc_hd__dfrtp_1
X_2431_ clknet_leaf_13_clk _0039_ net139 VGND VGND VDPWR VDPWR dig_ctrl_inst.cpu_inst.data\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_1313_ net154 net124 net78 VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.data_we\[12\]
+ sky130_fd_sc_hd__and3_2
X_1244_ _1002_ dig_ctrl_inst.spi_addr\[1\] VGND VGND VDPWR VDPWR _1092_ sky130_fd_sc_hd__or2_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[38\].gen_latches\[5\].p_latch net204 dig_ctrl_inst.latch_mem_inst.gclk\[38\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[38\]\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_47_76 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_8
X_2293_ _0751_ _0922_ _0920_ VGND VGND VDPWR VDPWR _0973_ sky130_fd_sc_hd__o21bai_1
X_2362_ dig_ctrl_inst.stb_dd _1039_ _0999_ VGND VGND VDPWR VDPWR _0989_ sky130_fd_sc_hd__a21o_1
XFILLER_0_74_333 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_97 VDPWR VGND VDPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_341 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_1175_ _1020_ _1022_ VGND VGND VDPWR VDPWR _1023_ sky130_fd_sc_hd__nand2_1
XANTENNA_12 dig_ctrl_inst.latch_mem_inst.gclk\[56\] VGND VGND VDPWR VDPWR sky130_fd_sc_hd__diode_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[27\].gen_latches\[3\].p_latch net217 dig_ctrl_inst.latch_mem_inst.gclk\[27\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[27\]\[3\] sky130_fd_sc_hd__dlxtp_1
XANTENNA_23 _0157_ VGND VGND VDPWR VDPWR sky130_fd_sc_hd__diode_2
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[11\].clock_buffer dig_ctrl_inst.latch_mem_inst.gen_gclk\[11\]._gclk
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.gclk\[11\] sky130_fd_sc_hd__clkbuf_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[16\].gen_latches\[1\].p_latch net232 dig_ctrl_inst.latch_mem_inst.gclk\[16\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[16\]\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_65_333 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_219 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_263 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_44_431 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[9\].gen_latches\[3\].p_latch net215 dig_ctrl_inst.latch_mem_inst.gclk\[9\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[9\]\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_17_57 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
Xinput10 ui_in[7] VGND VGND VDPWR VDPWR net10 sky130_fd_sc_hd__clkbuf_1
X_1862_ dig_ctrl_inst.latch_mem_inst.RAM\[30\]\[5\] net74 net69 _0159_ dig_ctrl_inst.latch_mem_inst.RAM\[62\]\[5\]
+ VGND VGND VDPWR VDPWR _0569_ sky130_fd_sc_hd__a32o_1
X_1931_ dig_ctrl_inst.latch_mem_inst.RAM\[1\]\[6\] net133 net124 net118 VGND VGND
+ VDPWR VDPWR _0637_ sky130_fd_sc_hd__and4_1
XFILLER_0_56_333 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_78 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_1793_ dig_ctrl_inst.latch_mem_inst.RAM\[39\]\[3\] _0139_ _0499_ _0500_ _0501_ VGND
+ VGND VDPWR VDPWR _0502_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_3_113 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XFILLER_0_58_75 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_42 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
X_2414_ clknet_leaf_13_clk _0022_ net141 VGND VGND VDPWR VDPWR dig_ctrl_inst.cpu_inst.ip\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_2345_ dig_ctrl_inst.cpu_inst.port_o\[0\] net390 _0987_ VGND VGND VDPWR VDPWR _0095_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_74_85 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_67_567 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1227_ dig_ctrl_inst.cpu_inst.ip\[0\] net293 _1030_ _1067_ _1074_ VGND VGND VDPWR
+ VDPWR _1075_ sky130_fd_sc_hd__a221oi_4
X_1158_ dig_ctrl_inst.cpu_inst.prev_state\[0\] VGND VGND VDPWR VDPWR _1007_ sky130_fd_sc_hd__inv_2
X_2276_ _0748_ _0956_ _0961_ _0955_ VGND VGND VDPWR VDPWR _0962_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_50_467 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_512 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_174 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_41_412 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_333 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_127 VDPWR VGND VDPWR VGND sky130_ef_sc_hd__decap_12
X_2061_ net257 net288 net261 VGND VGND VDPWR VDPWR _0754_ sky130_fd_sc_hd__or3b_4
XFILLER_0_28_56 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_2130_ _0257_ _0258_ _0821_ VGND VGND VDPWR VDPWR _0822_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_64_548 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_141 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
X_1914_ _0593_ _0598_ _0603_ _0620_ VGND VGND VDPWR VDPWR _0621_ sky130_fd_sc_hd__nor4_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[60\].gen_latches\[3\].p_latch net223 dig_ctrl_inst.latch_mem_inst.gclk\[60\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[60\]\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_71_111 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_1845_ dig_ctrl_inst.latch_mem_inst.RAM\[11\]\[4\] net124 net107 net92 VGND VGND
+ VDPWR VDPWR _0553_ sky130_fd_sc_hd__and4_1
X_1776_ dig_ctrl_inst.latch_mem_inst.RAM\[17\]\[3\] _0120_ _0482_ _0483_ _0484_ VGND
+ VGND VDPWR VDPWR _0485_ sky130_fd_sc_hd__a2111o_1
X_2328_ dig_ctrl_inst.spi_data_o\[0\] dig_ctrl_inst.spi_data_o\[1\] _0180_ VGND VGND
+ VDPWR VDPWR _0080_ sky130_fd_sc_hd__mux2_1
XFILLER_0_40_3 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_288 VDPWR VGND VDPWR VGND sky130_ef_sc_hd__decap_12
X_2259_ _0944_ _0945_ VGND VGND VDPWR VDPWR _0946_ sky130_fd_sc_hd__nand2_1
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[25\].clock_gate clknet_leaf_16_clk dig_ctrl_inst.latch_mem_inst.data_we\[25\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.gen_gclk\[25\]._gclk sky130_fd_sc_hd__dlclkp_1
XFILLER_0_50_306 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_260 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XFILLER_0_62_188 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_61_529 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_181 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1630_ dig_ctrl_inst.latch_mem_inst.RAM\[46\]\[1\] net72 net52 VGND VGND VDPWR VDPWR
+ _0341_ sky130_fd_sc_hd__and3_2
XFILLER_0_39_11 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
X_1492_ _0209_ dig_ctrl_inst.cpu_inst.ip\[1\] _0204_ VGND VGND VDPWR VDPWR _0020_
+ sky130_fd_sc_hd__mux2_1
X_1561_ net253 _0273_ VGND VGND VDPWR VDPWR _0274_ sky130_fd_sc_hd__xnor2_1
X_2113_ _0755_ _0805_ net165 _0754_ VGND VGND VDPWR VDPWR _0806_ sky130_fd_sc_hd__o2bb2a_1
X_2044_ net388 _0685_ _0741_ VGND VGND VDPWR VDPWR _0040_ sky130_fd_sc_hd__mux2_1
XFILLER_0_44_122 VDPWR VGND VDPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_141 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_188 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_8
X_1759_ dig_ctrl_inst.latch_mem_inst.RAM\[9\]\[3\] _1143_ _0158_ dig_ctrl_inst.latch_mem_inst.RAM\[61\]\[3\]
+ VGND VGND VDPWR VDPWR _0468_ sky130_fd_sc_hd__a22o_1
X_1828_ dig_ctrl_inst.latch_mem_inst.RAM\[45\]\[4\] net114 net80 net51 VGND VGND VDPWR
+ VDPWR _0536_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_9_218 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[53\].gen_latches\[2\].p_latch net226 dig_ctrl_inst.latch_mem_inst.gclk\[53\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[53\]\[2\] sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_0_162 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[42\].gen_latches\[0\].p_latch net243 dig_ctrl_inst.latch_mem_inst.gclk\[42\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[42\]\[0\] sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_74_610 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_57 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[30\].gen_latches\[7\].p_latch net187 dig_ctrl_inst.latch_mem_inst.gclk\[30\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[30\]\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_41_169 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_147 VDPWR VGND VDPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_136 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_1613_ dig_ctrl_inst.latch_mem_inst.RAM\[18\]\[0\] _0121_ _0151_ dig_ctrl_inst.latch_mem_inst.RAM\[53\]\[0\]
+ _0311_ VGND VGND VDPWR VDPWR _0325_ sky130_fd_sc_hd__a221o_1
XFILLER_0_26_188 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_244 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_1544_ _0254_ _0256_ VGND VGND VDPWR VDPWR _0257_ sky130_fd_sc_hd__nand2_1
XFILLER_0_14_306 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_317 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_339 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
X_1475_ dig_ctrl_inst.cpu_inst.r0\[4\] dig_ctrl_inst.cpu_inst.port_o\[4\] _0176_ VGND
+ VGND VDPWR VDPWR _0015_ sky130_fd_sc_hd__mux2_1
Xfanout219 net329 VGND VGND VDPWR VDPWR net219 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_5_78 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
Xfanout208 net209 VGND VGND VDPWR VDPWR net208 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_37_389 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2027_ dig_ctrl_inst.latch_mem_inst.RAM\[21\]\[7\] _0124_ _0150_ dig_ctrl_inst.latch_mem_inst.RAM\[52\]\[7\]
+ VGND VGND VDPWR VDPWR _0732_ sky130_fd_sc_hd__a22o_1
XFILLER_0_64_239 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_147 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_17_Left_95 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_144 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[57\].gen_latches\[3\].p_latch net220 dig_ctrl_inst.latch_mem_inst.gclk\[57\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[57\]\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_20_309 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_28_334 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[46\].gen_latches\[1\].p_latch net234 dig_ctrl_inst.latch_mem_inst.gclk\[46\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[46\]\[1\] sky130_fd_sc_hd__dlxtp_1
Xinput8 ui_in[5] VGND VGND VDPWR VDPWR net8 sky130_fd_sc_hd__clkbuf_1
X_1260_ net267 dig_ctrl_inst.cpu_inst.r2\[5\] VGND VGND VDPWR VDPWR _1108_ sky130_fd_sc_hd__and2b_1
X_1191_ net248 dig_ctrl_inst.cpu_inst.cpu_state\[1\] _0999_ VGND VGND VDPWR VDPWR
+ _1039_ sky130_fd_sc_hd__nor3_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[1\].gen_latches\[5\].p_latch net202 dig_ctrl_inst.latch_mem_inst.gclk\[1\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[1\]\[5\] sky130_fd_sc_hd__dlxtp_1
X_1527_ _0238_ _0239_ VGND VGND VDPWR VDPWR _0240_ sky130_fd_sc_hd__or2_1
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[4\].clock_gate clknet_leaf_19_clk dig_ctrl_inst.latch_mem_inst.data_we\[4\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.gen_gclk\[4\]._gclk sky130_fd_sc_hd__dlclkp_1
X_1458_ _1096_ _0189_ _0188_ _0184_ VGND VGND VDPWR VDPWR _0006_ sky130_fd_sc_hd__o211a_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[23\].gen_latches\[6\].p_latch net192 dig_ctrl_inst.latch_mem_inst.gclk\[23\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[23\]\[6\] sky130_fd_sc_hd__dlxtp_1
X_1389_ net96 net43 VGND VGND VDPWR VDPWR _0150_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_25_315 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[12\].gen_latches\[4\].p_latch net214 dig_ctrl_inst.latch_mem_inst.gclk\[12\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[12\]\[4\] sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[39\].gen_latches\[0\].p_latch net245 dig_ctrl_inst.latch_mem_inst.gclk\[39\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[39\]\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_22_36 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
X_2361_ dig_ctrl_inst.cpu_inst.port_o\[7\] net353 _0988_ VGND VGND VDPWR VDPWR _0110_
+ sky130_fd_sc_hd__mux2_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[5\].gen_latches\[6\].p_latch net198 dig_ctrl_inst.latch_mem_inst.gclk\[5\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[5\]\[6\] sky130_fd_sc_hd__dlxtp_1
X_2430_ clknet_leaf_13_clk _0038_ net139 VGND VGND VDPWR VDPWR dig_ctrl_inst.cpu_inst.data\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_1312_ net125 net79 VGND VGND VDPWR VDPWR _1148_ sky130_fd_sc_hd__and2_1
X_2292_ net359 _0972_ _0967_ VGND VGND VDPWR VDPWR _0057_ sky130_fd_sc_hd__mux2_1
X_1243_ _1039_ net162 VGND VGND VDPWR VDPWR _1091_ sky130_fd_sc_hd__and2_1
XFILLER_0_47_99 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_1174_ net264 net265 VGND VGND VDPWR VDPWR _1022_ sky130_fd_sc_hd__and2b_1
XFILLER_0_63_76 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XANTENNA_13 dig_ctrl_inst.latch_mem_inst.gclk\[56\] VGND VGND VDPWR VDPWR sky130_fd_sc_hd__diode_2
XFILLER_0_2_79 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[50\].clock_buffer dig_ctrl_inst.latch_mem_inst.gen_gclk\[50\]._gclk
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.gclk\[50\] sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_25_Left_103 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XFILLER_0_70_3 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
XANTENNA_24 _0157_ VGND VGND VDPWR VDPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_166 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_8
Xdig_ctrl_inst.latch_mem_inst.gen_words\[27\].gen_latches\[7\].p_latch net189 dig_ctrl_inst.latch_mem_inst.gclk\[27\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[27\]\[7\] sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_34_Left_112 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_43_Left_121 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[16\].gen_latches\[5\].p_latch net199 dig_ctrl_inst.latch_mem_inst.gclk\[16\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[16\]\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_18_250 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_52_Left_130 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[32\].clock_gate clknet_leaf_15_clk dig_ctrl_inst.latch_mem_inst.data_we\[32\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.gen_gclk\[32\]._gclk sky130_fd_sc_hd__dlclkp_1
XFILLER_0_0_309 VDPWR VGND VDPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_57 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_35 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_1930_ dig_ctrl_inst.latch_mem_inst.RAM\[16\]\[6\] net128 net62 VGND VGND VDPWR VDPWR
+ _0636_ sky130_fd_sc_hd__and3_2
Xinput11 uio_in[0] VGND VGND VDPWR VDPWR net11 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_71_337 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_1861_ dig_ctrl_inst.latch_mem_inst.RAM\[11\]\[5\] _1145_ _0155_ dig_ctrl_inst.latch_mem_inst.RAM\[58\]\[5\]
+ _0567_ VGND VGND VDPWR VDPWR _0568_ sky130_fd_sc_hd__a221o_1
X_1792_ dig_ctrl_inst.latch_mem_inst.RAM\[56\]\[3\] net87 net46 VGND VGND VDPWR VDPWR
+ _0501_ sky130_fd_sc_hd__and3_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[9\].gen_latches\[7\].p_latch net183 dig_ctrl_inst.latch_mem_inst.gclk\[9\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[9\]\[7\] sky130_fd_sc_hd__dlxtp_1
X_2344_ dig_ctrl_inst.cpu_inst.port_stb_o _0802_ VGND VGND VDPWR VDPWR _0987_ sky130_fd_sc_hd__nand2_4
X_2413_ clknet_leaf_9_clk _0021_ net141 VGND VGND VDPWR VDPWR dig_ctrl_inst.cpu_inst.ip\[2\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_1_0__f_clk clknet_0_clk VGND VGND VDPWR VDPWR clknet_1_0__leaf_clk sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_67_568 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1226_ _1039_ net165 net249 VGND VGND VDPWR VDPWR _1074_ sky130_fd_sc_hd__a21o_1
X_1157_ dig_ctrl_inst.cpu_inst.ip\[5\] VGND VGND VDPWR VDPWR _1006_ sky130_fd_sc_hd__inv_2
X_2275_ _0749_ _0956_ _0960_ VGND VGND VDPWR VDPWR _0961_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_15_275 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_297 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_513 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_413 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_337 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
XFILLER_0_53_304 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_24 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_5_Left_83 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_139 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_64_549 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_23 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
X_2060_ net257 net287 net261 VGND VGND VDPWR VDPWR _0753_ sky130_fd_sc_hd__nor3b_1
X_1913_ _0607_ _0611_ _0615_ _0619_ VGND VGND VDPWR VDPWR _0620_ sky130_fd_sc_hd__or4_1
X_1844_ dig_ctrl_inst.latch_mem_inst.RAM\[12\]\[4\] net124 net78 VGND VGND VDPWR VDPWR
+ _0552_ sky130_fd_sc_hd__and3_2
X_1775_ dig_ctrl_inst.latch_mem_inst.RAM\[49\]\[3\] net133 net117 net46 VGND VGND
+ VDPWR VDPWR _0484_ sky130_fd_sc_hd__and4_1
XFILLER_0_12_223 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[60\].gen_latches\[7\].p_latch net188 dig_ctrl_inst.latch_mem_inst.gclk\[60\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[60\]\[7\] sky130_fd_sc_hd__dlxtp_1
X_2327_ net345 dig_ctrl_inst.spi_data_o\[0\] _0180_ VGND VGND VDPWR VDPWR _0079_ sky130_fd_sc_hd__mux2_1
X_2258_ _0227_ _0921_ VGND VGND VDPWR VDPWR _0945_ sky130_fd_sc_hd__or2_1
XFILLER_0_33_3 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
X_1209_ net268 dig_ctrl_inst.cpu_inst.r2\[2\] VGND VGND VDPWR VDPWR _1057_ sky130_fd_sc_hd__and2b_1
X_2189_ net166 net165 net162 _1045_ VGND VGND VDPWR VDPWR _0879_ sky130_fd_sc_hd__a31o_1
XFILLER_0_7_294 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_3_182 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_131 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_8
X_1560_ _0268_ _0272_ _0262_ VGND VGND VDPWR VDPWR _0273_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_77_630 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2112_ dig_ctrl_inst.synchronizer_port_i_inst\[0\].out _0802_ _0804_ dig_ctrl_inst.spi_data_o\[0\]
+ _0803_ VGND VGND VDPWR VDPWR _0805_ sky130_fd_sc_hd__a221o_1
X_1491_ _0207_ _0208_ _0174_ VGND VGND VDPWR VDPWR _0209_ sky130_fd_sc_hd__mux2_1
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[43\].clock_buffer dig_ctrl_inst.latch_mem_inst.gen_gclk\[43\]._gclk
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.gclk\[43\] sky130_fd_sc_hd__clkbuf_4
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[9\].clock_gate clknet_leaf_15_clk dig_ctrl_inst.latch_mem_inst.data_we\[9\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.gen_gclk\[9\]._gclk sky130_fd_sc_hd__dlclkp_1
X_2043_ dig_ctrl_inst.cpu_inst.data\[5\] _0622_ _0741_ VGND VGND VDPWR VDPWR _0039_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_44_134 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_197 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
X_1827_ dig_ctrl_inst.latch_mem_inst.RAM\[61\]\[4\] net114 net80 net42 VGND VGND VDPWR
+ VDPWR _0535_ sky130_fd_sc_hd__and4_1
XFILLER_0_17_337 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
X_1689_ dig_ctrl_inst.latch_mem_inst.RAM\[62\]\[2\] net74 net49 VGND VGND VDPWR VDPWR
+ _0399_ sky130_fd_sc_hd__and3_2
XTAP_TAPCELL_ROW_9_219 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1758_ dig_ctrl_inst.latch_mem_inst.RAM\[52\]\[3\] _0150_ _0152_ dig_ctrl_inst.latch_mem_inst.RAM\[54\]\[3\]
+ VGND VGND VDPWR VDPWR _0467_ sky130_fd_sc_hd__a22o_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[53\].gen_latches\[6\].p_latch net194 dig_ctrl_inst.latch_mem_inst.gclk\[53\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[53\]\[6\] sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_0_163 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[42\].gen_latches\[4\].p_latch net214 dig_ctrl_inst.latch_mem_inst.gclk\[42\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[42\]\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_50_126 VDPWR VGND VDPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_611 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[31\].gen_latches\[2\].p_latch net225 dig_ctrl_inst.latch_mem_inst.gclk\[31\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[31\]\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_41_57 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_112 VDPWR VGND VDPWR VGND sky130_ef_sc_hd__decap_12
X_1474_ dig_ctrl_inst.cpu_inst.r0\[3\] dig_ctrl_inst.cpu_inst.port_o\[3\] _0176_ VGND
+ VGND VDPWR VDPWR _0014_ sky130_fd_sc_hd__mux2_1
X_1612_ _0306_ _0308_ _0322_ _0323_ VGND VGND VDPWR VDPWR _0324_ sky130_fd_sc_hd__or4_1
XFILLER_0_41_159 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[20\].gen_latches\[0\].p_latch net245 dig_ctrl_inst.latch_mem_inst.gclk\[20\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[20\]\[0\] sky130_fd_sc_hd__dlxtp_1
Xfanout209 net323 VGND VGND VDPWR VDPWR net209 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_1_289 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_223 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_1543_ net163 net161 VGND VGND VDPWR VDPWR _0256_ sky130_fd_sc_hd__or2_1
XFILLER_0_5_57 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_323 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
X_2026_ dig_ctrl_inst.latch_mem_inst.RAM\[23\]\[7\] _0126_ _0688_ _0689_ _0704_ VGND
+ VGND VDPWR VDPWR _0731_ sky130_fd_sc_hd__a2111o_1
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[37\].clock_gate clknet_leaf_19_clk dig_ctrl_inst.latch_mem_inst.data_we\[37\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.gen_gclk\[37\]._gclk sky130_fd_sc_hd__dlclkp_1
XFILLER_0_32_137 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_189 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[57\].gen_latches\[7\].p_latch net186 dig_ctrl_inst.latch_mem_inst.gclk\[57\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[57\]\[7\] sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_28_335 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_262 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[2\].gen_latches\[0\].p_latch net245 dig_ctrl_inst.latch_mem_inst.gclk\[2\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[2\]\[0\] sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[46\].gen_latches\[5\].p_latch net201 dig_ctrl_inst.latch_mem_inst.gclk\[46\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[46\]\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_31_181 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
Xinput9 ui_in[6] VGND VGND VDPWR VDPWR net9 sky130_fd_sc_hd__clkbuf_1
X_1190_ _1010_ _1025_ _1036_ VGND VGND VDPWR VDPWR _1038_ sky130_fd_sc_hd__and3_2
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[0\].clock_buffer dig_ctrl_inst.latch_mem_inst.gen_gclk\[0\]._gclk
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.gclk\[0\] sky130_fd_sc_hd__clkbuf_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[35\].gen_latches\[3\].p_latch net216 dig_ctrl_inst.latch_mem_inst.gclk\[35\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[35\]\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_52_78 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_262 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[24\].gen_latches\[1\].p_latch net233 dig_ctrl_inst.latch_mem_inst.gclk\[24\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[24\]\[1\] sky130_fd_sc_hd__dlxtp_1
X_1457_ dig_ctrl_inst.spi_addr\[0\] dig_ctrl_inst.spi_addr\[1\] VGND VGND VDPWR VDPWR
+ _0189_ sky130_fd_sc_hd__nand2_1
X_1526_ _1118_ net159 VGND VGND VDPWR VDPWR _0239_ sky130_fd_sc_hd__nor2_1
X_1388_ net150 _0149_ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.data_we\[51\]
+ sky130_fd_sc_hd__and2_1
X_2009_ dig_ctrl_inst.latch_mem_inst.RAM\[31\]\[7\] _0132_ _0277_ dig_ctrl_inst.latch_mem_inst.RAM\[4\]\[7\]
+ VGND VGND VDPWR VDPWR _0714_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_33_360 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_316 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_321 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[6\].gen_latches\[1\].p_latch net232 dig_ctrl_inst.latch_mem_inst.gclk\[6\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[6\]\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_36_295 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_2360_ dig_ctrl_inst.cpu_inst.port_o\[6\] net383 _0988_ VGND VGND VDPWR VDPWR _0109_
+ sky130_fd_sc_hd__mux2_1
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[36\].clock_buffer dig_ctrl_inst.latch_mem_inst.gen_gclk\[36\]._gclk
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.gclk\[36\] sky130_fd_sc_hd__clkbuf_4
X_1311_ _1075_ _1077_ net134 net135 _1047_ VGND VGND VDPWR VDPWR _1147_ sky130_fd_sc_hd__o2111a_1
X_2291_ _0751_ _0903_ _0900_ VGND VGND VDPWR VDPWR _0972_ sky130_fd_sc_hd__o21ai_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[39\].gen_latches\[4\].p_latch net213 dig_ctrl_inst.latch_mem_inst.gclk\[39\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[39\]\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_63_44 VDPWR VGND VDPWR VGND sky130_ef_sc_hd__decap_12
X_1173_ net267 net263 VGND VGND VDPWR VDPWR _1021_ sky130_fd_sc_hd__nor2_4
X_1242_ net181 _1086_ _1087_ _1088_ _1089_ VGND VGND VDPWR VDPWR _1090_ sky130_fd_sc_hd__o41a_1
XPHY_EDGE_ROW_10_Right_10 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[28\].gen_latches\[2\].p_latch net230 dig_ctrl_inst.latch_mem_inst.gclk\[28\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[28\]\[2\] sky130_fd_sc_hd__dlxtp_1
XANTENNA_25 _0187_ VGND VGND VDPWR VDPWR sky130_fd_sc_hd__diode_2
XANTENNA_14 dig_ctrl_inst.latch_mem_inst.gclk\[6\] VGND VGND VDPWR VDPWR sky130_fd_sc_hd__diode_2
XFILLER_0_63_3 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_232 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_2489_ clknet_leaf_4_clk _0088_ net177 VGND VGND VDPWR VDPWR dig_ctrl_inst.spi_data_i\[1\]
+ sky130_fd_sc_hd__dfrtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[17\].gen_latches\[0\].p_latch net243 dig_ctrl_inst.latch_mem_inst.gclk\[17\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[17\]\[0\] sky130_fd_sc_hd__dlxtp_1
X_1509_ net160 dig_ctrl_inst.cpu_inst.data\[5\] _0198_ VGND VGND VDPWR VDPWR _0223_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_313 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_1860_ dig_ctrl_inst.latch_mem_inst.RAM\[25\]\[5\] _0128_ _0153_ dig_ctrl_inst.latch_mem_inst.RAM\[55\]\[5\]
+ VGND VGND VDPWR VDPWR _0567_ sky130_fd_sc_hd__a22o_1
Xinput12 uio_in[1] VGND VGND VDPWR VDPWR net12 sky130_fd_sc_hd__clkbuf_1
X_1791_ dig_ctrl_inst.latch_mem_inst.RAM\[36\]\[3\] net98 net56 VGND VGND VDPWR VDPWR
+ _0500_ sky130_fd_sc_hd__and3_2
X_2343_ dig_ctrl_inst.cpu_inst.port_o\[7\] net351 _0986_ VGND VGND VDPWR VDPWR _0094_
+ sky130_fd_sc_hd__mux2_1
X_2412_ clknet_leaf_9_clk _0020_ net141 VGND VGND VDPWR VDPWR dig_ctrl_inst.cpu_inst.ip\[1\]
+ sky130_fd_sc_hd__dfrtp_2
X_2274_ _0172_ _0233_ _0792_ _0959_ VGND VGND VDPWR VDPWR _0960_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_67_569 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1225_ net181 _1071_ _1070_ _1069_ _1072_ VGND VGND VDPWR VDPWR _1073_ sky130_fd_sc_hd__o41a_1
Xclkbuf_leaf_17_clk clknet_1_0__leaf_clk VGND VGND VDPWR VDPWR clknet_leaf_17_clk
+ sky130_fd_sc_hd__clkbuf_8
X_1156_ dig_ctrl_inst.cpu_inst.ip\[4\] VGND VGND VDPWR VDPWR _1005_ sky130_fd_sc_hd__inv_2
XFILLER_0_62_338 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
XFILLER_0_59_195 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_184 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_1989_ dig_ctrl_inst.latch_mem_inst.RAM\[38\]\[7\] net93 net51 VGND VGND VDPWR VDPWR
+ _0694_ sky130_fd_sc_hd__and3_2
XFILLER_0_15_210 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_58_514 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_313 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_202 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_69 VDPWR VGND VDPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_279 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_72_594 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_56 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_34 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_6
X_1843_ _0538_ _0542_ _0546_ _0550_ VGND VGND VDPWR VDPWR _0551_ sky130_fd_sc_hd__or4_1
XFILLER_0_29_335 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_1912_ dig_ctrl_inst.latch_mem_inst.RAM\[9\]\[5\] _1143_ _0616_ _0617_ _0618_ VGND
+ VGND VDPWR VDPWR _0619_ sky130_fd_sc_hd__a2111o_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[61\].gen_latches\[2\].p_latch net224 dig_ctrl_inst.latch_mem_inst.gclk\[61\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[61\]\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_69_43 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_6_clk clknet_1_1__leaf_clk VGND VGND VDPWR VDPWR clknet_leaf_6_clk sky130_fd_sc_hd__clkbuf_8
X_1774_ dig_ctrl_inst.latch_mem_inst.RAM\[45\]\[3\] net117 net81 net56 VGND VGND VDPWR
+ VDPWR _0483_ sky130_fd_sc_hd__and4_1
XPHY_EDGE_ROW_71_Left_149 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
X_2326_ net174 dig_ctrl_inst.spi_receiver_inst.spi_cnt\[2\] _0182_ _0985_ VGND VGND
+ VDPWR VDPWR _0078_ sky130_fd_sc_hd__a31o_1
X_1208_ net268 net263 dig_ctrl_inst.cpu_inst.r3\[2\] VGND VGND VDPWR VDPWR _1056_
+ sky130_fd_sc_hd__and3_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[50\].gen_latches\[0\].p_latch net246 dig_ctrl_inst.latch_mem_inst.gclk\[50\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[50\]\[0\] sky130_fd_sc_hd__dlxtp_1
X_2257_ net138 _0921_ VGND VGND VDPWR VDPWR _0944_ sky130_fd_sc_hd__nand2_1
XFILLER_0_26_3 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
X_2188_ _1045_ net166 net165 net162 VGND VGND VDPWR VDPWR _0878_ sky130_fd_sc_hd__and4_1
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[44\].clock_gate clknet_leaf_19_clk dig_ctrl_inst.latch_mem_inst.data_we\[44\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.gen_gclk\[44\]._gclk sky130_fd_sc_hd__dlclkp_1
XTAP_TAPCELL_ROW_3_183 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_113 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
XFILLER_0_53_124 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
XFILLER_0_38_187 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[29\].clock_buffer dig_ctrl_inst.latch_mem_inst.gen_gclk\[29\]._gclk
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.gclk\[29\] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_39_57 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
X_1490_ dig_ctrl_inst.cpu_inst.ip\[0\] dig_ctrl_inst.cpu_inst.ip\[1\] VGND VGND VDPWR
+ VDPWR _0208_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_77_631 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2111_ _0799_ dig_ctrl_inst.cpu_inst.data\[0\] dig_ctrl_inst.cpu_inst.data\[1\] _0801_
+ VGND VGND VDPWR VDPWR _0804_ sky130_fd_sc_hd__and4bb_4
X_2042_ dig_ctrl_inst.cpu_inst.data\[4\] _0565_ _0741_ VGND VGND VDPWR VDPWR _0038_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_71_88 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_66 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_55 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_8_Right_8 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
X_1826_ _0523_ _0527_ _0529_ _0533_ VGND VGND VDPWR VDPWR _0534_ sky130_fd_sc_hd__or4_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[54\].gen_latches\[1\].p_latch net237 dig_ctrl_inst.latch_mem_inst.gclk\[54\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[54\]\[1\] sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_39_Right_39 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_341 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_1688_ net263 _0398_ _0276_ VGND VGND VDPWR VDPWR _0027_ sky130_fd_sc_hd__mux2_1
X_1757_ dig_ctrl_inst.latch_mem_inst.RAM\[25\]\[3\] _0128_ _0151_ dig_ctrl_inst.latch_mem_inst.RAM\[53\]\[3\]
+ _0465_ VGND VGND VDPWR VDPWR _0466_ sky130_fd_sc_hd__a221o_1
X_2309_ net360 _0968_ _0977_ VGND VGND VDPWR VDPWR _0069_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_48_Right_48 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_91 VDPWR VGND VDPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_164 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_57_Right_57 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_138 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_116 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_341 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_66_Right_66 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
X_1611_ dig_ctrl_inst.latch_mem_inst.RAM\[11\]\[0\] _1145_ _0117_ dig_ctrl_inst.latch_mem_inst.RAM\[15\]\[0\]
+ _0309_ VGND VGND VDPWR VDPWR _0323_ sky130_fd_sc_hd__a221o_1
XFILLER_0_26_124 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[31\].gen_latches\[6\].p_latch net191 dig_ctrl_inst.latch_mem_inst.gclk\[31\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[31\]\[6\] sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_75_Right_75 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
X_1473_ dig_ctrl_inst.cpu_inst.r0\[2\] dig_ctrl_inst.cpu_inst.port_o\[2\] _0176_ VGND
+ VGND VDPWR VDPWR _0013_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_279 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_1542_ net163 net161 VGND VGND VDPWR VDPWR _0255_ sky130_fd_sc_hd__nor2_1
XFILLER_0_66_66 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[20\].gen_latches\[4\].p_latch net212 dig_ctrl_inst.latch_mem_inst.gclk\[20\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[20\]\[4\] sky130_fd_sc_hd__dlxtp_1
X_2025_ dig_ctrl_inst.latch_mem_inst.RAM\[9\]\[7\] _1143_ _0135_ dig_ctrl_inst.latch_mem_inst.RAM\[33\]\[7\]
+ _0699_ VGND VGND VDPWR VDPWR _0730_ sky130_fd_sc_hd__a221o_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[58\].gen_latches\[2\].p_latch net229 dig_ctrl_inst.latch_mem_inst.gclk\[58\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[58\]\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_9_313 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_335 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_70 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_1809_ dig_ctrl_inst.latch_mem_inst.RAM\[7\]\[4\] _1139_ _0514_ _0515_ _0516_ VGND
+ VGND VDPWR VDPWR _0517_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_13_341 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[47\].gen_latches\[0\].p_latch net242 dig_ctrl_inst.latch_mem_inst.gclk\[47\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[47\]\[0\] sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_36_380 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[2\].gen_latches\[4\].p_latch net210 dig_ctrl_inst.latch_mem_inst.gclk\[2\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[2\]\[4\] sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[35\].gen_latches\[7\].p_latch net184 dig_ctrl_inst.latch_mem_inst.gclk\[35\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[35\]\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_6_305 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[24\].gen_latches\[5\].p_latch net203 dig_ctrl_inst.latch_mem_inst.gclk\[24\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[24\]\[5\] sky130_fd_sc_hd__dlxtp_1
X_1456_ dig_ctrl_inst.spi_addr\[0\] _0185_ dig_ctrl_inst.spi_addr\[1\] VGND VGND VDPWR
+ VDPWR _0188_ sky130_fd_sc_hd__a21o_1
X_1525_ _1118_ net159 VGND VGND VDPWR VDPWR _0238_ sky130_fd_sc_hd__and2_1
X_1387_ net131 net102 net43 VGND VGND VDPWR VDPWR _0149_ sky130_fd_sc_hd__and3_2
X_2008_ dig_ctrl_inst.latch_mem_inst.RAM\[20\]\[7\] _0123_ _0136_ dig_ctrl_inst.latch_mem_inst.RAM\[34\]\[7\]
+ VGND VGND VDPWR VDPWR _0713_ sky130_fd_sc_hd__a22o_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[13\].gen_latches\[3\].p_latch net217 dig_ctrl_inst.latch_mem_inst.gclk\[13\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[13\]\[3\] sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_25_317 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_361 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_165 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[6\].gen_latches\[5\].p_latch net204 dig_ctrl_inst.latch_mem_inst.gclk\[6\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[6\]\[5\] sky130_fd_sc_hd__dlxtp_1
X_1310_ _1047_ net135 VGND VGND VDPWR VDPWR _1146_ sky130_fd_sc_hd__and2_4
X_2290_ net375 _0971_ _0967_ VGND VGND VDPWR VDPWR _0056_ sky130_fd_sc_hd__mux2_1
X_1241_ net266 net262 dig_ctrl_inst.cpu_inst.r0\[1\] VGND VGND VDPWR VDPWR _1089_
+ sky130_fd_sc_hd__or3_1
X_1172_ net286 _1019_ VGND VGND VDPWR VDPWR _1020_ sky130_fd_sc_hd__nor2_1
XFILLER_0_2_15 VDPWR VGND VDPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_26 _1039_ VGND VGND VDPWR VDPWR sky130_fd_sc_hd__diode_2
XANTENNA_15 dig_ctrl_inst.spi_data_i\[1\] VGND VGND VDPWR VDPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_342 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[28\].gen_latches\[6\].p_latch net194 dig_ctrl_inst.latch_mem_inst.gclk\[28\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[28\]\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_6_102 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_3 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_141 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_2488_ clknet_leaf_5_clk _0087_ net177 VGND VGND VDPWR VDPWR dig_ctrl_inst.spi_data_i\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_1439_ _0176_ VGND VGND VDPWR VDPWR _0000_ sky130_fd_sc_hd__inv_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[17\].gen_latches\[4\].p_latch net211 dig_ctrl_inst.latch_mem_inst.gclk\[17\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[17\]\[4\] sky130_fd_sc_hd__dlxtp_1
X_1508_ _0222_ _0204_ dig_ctrl_inst.cpu_inst.ip\[4\] _0220_ VGND VGND VDPWR VDPWR
+ _0023_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_65_303 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[49\].clock_gate clknet_leaf_19_clk dig_ctrl_inst.latch_mem_inst.data_we\[49\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.gen_gclk\[49\]._gclk sky130_fd_sc_hd__dlclkp_1
Xinput13 uio_in[3] VGND VGND VDPWR VDPWR net13 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_71_306 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_141 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
X_1790_ dig_ctrl_inst.latch_mem_inst.RAM\[37\]\[3\] net117 net100 net56 VGND VGND
+ VDPWR VDPWR _0499_ sky130_fd_sc_hd__and4_1
X_2411_ clknet_leaf_13_clk _0019_ net139 VGND VGND VDPWR VDPWR dig_ctrl_inst.cpu_inst.ip\[0\]
+ sky130_fd_sc_hd__dfrtp_4
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[51\].clock_gate clknet_leaf_13_clk dig_ctrl_inst.latch_mem_inst.data_we\[51\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.gen_gclk\[51\]._gclk sky130_fd_sc_hd__dlclkp_1
X_2342_ dig_ctrl_inst.cpu_inst.port_o\[6\] net350 _0986_ VGND VGND VDPWR VDPWR _0093_
+ sky130_fd_sc_hd__mux2_1
X_1224_ dig_ctrl_inst.cpu_inst.r0\[0\] net265 net262 VGND VGND VDPWR VDPWR _1072_
+ sky130_fd_sc_hd__or3_1
X_2273_ dig_ctrl_inst.cpu_inst.data\[7\] _0743_ _0825_ net138 _0958_ VGND VGND VDPWR
+ VDPWR _0959_ sky130_fd_sc_hd__a221o_1
XFILLER_0_74_99 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_1155_ dig_ctrl_inst.cpu_inst.ip\[3\] VGND VGND VDPWR VDPWR _1004_ sky130_fd_sc_hd__inv_2
XFILLER_0_62_306 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
X_1988_ dig_ctrl_inst.latch_mem_inst.RAM\[53\]\[7\] net114 net99 net42 VGND VGND VDPWR
+ VDPWR _0693_ sky130_fd_sc_hd__and4_1
XFILLER_0_2_160 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_515 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_188 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
Xfanout190 net328 VGND VGND VDPWR VDPWR net190 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_28_48 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_72_595 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1842_ dig_ctrl_inst.latch_mem_inst.RAM\[5\]\[4\] _0278_ _0547_ _0548_ _0549_ VGND
+ VGND VDPWR VDPWR _0550_ sky130_fd_sc_hd__a2111o_1
X_1773_ dig_ctrl_inst.latch_mem_inst.RAM\[27\]\[3\] net104 net91 net66 VGND VGND VDPWR
+ VDPWR _0482_ sky130_fd_sc_hd__and4_1
X_1911_ dig_ctrl_inst.latch_mem_inst.RAM\[45\]\[5\] net115 net80 net52 VGND VGND VDPWR
+ VDPWR _0618_ sky130_fd_sc_hd__and4_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[61\].gen_latches\[6\].p_latch net191 dig_ctrl_inst.latch_mem_inst.gclk\[61\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[61\]\[6\] sky130_fd_sc_hd__dlxtp_1
X_2325_ net174 dig_ctrl_inst.spi_receiver_inst.stb_o VGND VGND VDPWR VDPWR _0985_
+ sky130_fd_sc_hd__and2b_1
X_1207_ _1010_ _1025_ _1054_ VGND VGND VDPWR VDPWR _1055_ sky130_fd_sc_hd__and3_2
X_2187_ _0866_ _0876_ VGND VGND VDPWR VDPWR _0877_ sky130_fd_sc_hd__and2_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[50\].gen_latches\[4\].p_latch net210 dig_ctrl_inst.latch_mem_inst.gclk\[50\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[50\]\[4\] sky130_fd_sc_hd__dlxtp_1
X_2256_ _0788_ _0928_ _0932_ _0942_ VGND VGND VDPWR VDPWR _0943_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_63_540 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_133 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_3_184 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_169 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_27 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_339 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_77_632 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2110_ dig_ctrl_inst.cpu_inst.data\[0\] dig_ctrl_inst.port_ms_sync_i _0800_ _0801_
+ VGND VGND VDPWR VDPWR _0803_ sky130_fd_sc_hd__and4_1
XFILLER_0_55_57 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_46 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_2041_ dig_ctrl_inst.cpu_inst.data\[3\] _0505_ _0741_ VGND VGND VDPWR VDPWR _0037_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_17_264 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_147 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_309 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_1756_ dig_ctrl_inst.latch_mem_inst.RAM\[40\]\[3\] net86 net53 VGND VGND VDPWR VDPWR
+ _0465_ sky130_fd_sc_hd__and3_2
X_1825_ dig_ctrl_inst.latch_mem_inst.RAM\[25\]\[4\] _0128_ _0530_ _0531_ _0532_ VGND
+ VGND VDPWR VDPWR _0533_ sky130_fd_sc_hd__a2111o_1
X_1687_ dig_ctrl_inst.latch_mem_inst.RAM\[0\]\[1\] _0288_ _0384_ _0397_ VGND VGND
+ VDPWR VDPWR _0398_ sky130_fd_sc_hd__o22a_1
X_2308_ net265 net264 _0175_ _0756_ VGND VGND VDPWR VDPWR _0977_ sky130_fd_sc_hd__and4_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[54\].gen_latches\[5\].p_latch net202 dig_ctrl_inst.latch_mem_inst.gclk\[54\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[54\]\[5\] sky130_fd_sc_hd__dlxtp_1
X_2239_ dig_ctrl_inst.cpu_inst.r0\[6\] net41 VGND VGND VDPWR VDPWR _0926_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_0_165 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_169 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_6
Xdig_ctrl_inst.latch_mem_inst.gen_words\[43\].gen_latches\[3\].p_latch net218 dig_ctrl_inst.latch_mem_inst.gclk\[43\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[43\]\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_23_309 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_3 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_8_210 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_90 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[32\].gen_latches\[1\].p_latch net233 dig_ctrl_inst.latch_mem_inst.gclk\[32\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[32\]\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_58_228 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_1610_ _0310_ _0321_ VGND VGND VDPWR VDPWR _0322_ sky130_fd_sc_hd__or2_1
X_1472_ dig_ctrl_inst.cpu_inst.r0\[1\] dig_ctrl_inst.cpu_inst.port_o\[1\] _0176_ VGND
+ VGND VDPWR VDPWR _0012_ sky130_fd_sc_hd__mux2_1
X_1541_ net163 net161 VGND VGND VDPWR VDPWR _0254_ sky130_fd_sc_hd__nand2_1
X_2024_ _0717_ _0722_ _0724_ VGND VGND VDPWR VDPWR _0729_ sky130_fd_sc_hd__or3_1
XFILLER_0_17_169 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_1808_ dig_ctrl_inst.latch_mem_inst.RAM\[27\]\[4\] net108 _1140_ net68 VGND VGND
+ VDPWR VDPWR _0516_ sky130_fd_sc_hd__and4_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[58\].gen_latches\[6\].p_latch net198 dig_ctrl_inst.latch_mem_inst.gclk\[58\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[58\]\[6\] sky130_fd_sc_hd__dlxtp_1
X_1739_ _0434_ _0435_ _0448_ _0288_ dig_ctrl_inst.latch_mem_inst.RAM\[0\]\[2\] VGND
+ VGND VDPWR VDPWR _0449_ sky130_fd_sc_hd__o32a_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[47\].gen_latches\[4\].p_latch net211 dig_ctrl_inst.latch_mem_inst.gclk\[47\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[47\]\[4\] sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_36_381 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_275 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[56\].clock_gate clknet_leaf_0_clk dig_ctrl_inst.latch_mem_inst.data_we\[56\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.gen_gclk\[56\]._gclk sky130_fd_sc_hd__dlclkp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[36\].gen_latches\[2\].p_latch net226 dig_ctrl_inst.latch_mem_inst.gclk\[36\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[36\]\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_36_59 VDPWR VGND VDPWR VGND sky130_ef_sc_hd__decap_12
Xdig_ctrl_inst.latch_mem_inst.gen_words\[25\].gen_latches\[0\].p_latch net240 dig_ctrl_inst.latch_mem_inst.gclk\[25\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[25\]\[0\] sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_input_latches\[0\].n_latch dig_ctrl_inst.data_out\[0\]
+ clknet_leaf_2_clk VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.wdata\[0\]
+ sky130_fd_sc_hd__dlxtn_1
XFILLER_0_54_231 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_33 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_1524_ _0230_ _0236_ VGND VGND VDPWR VDPWR _0237_ sky130_fd_sc_hd__nand2_1
XFILLER_0_22_172 VDPWR VGND VDPWR VGND sky130_ef_sc_hd__decap_12
X_1455_ net382 _0185_ _0187_ VGND VGND VDPWR VDPWR _0005_ sky130_fd_sc_hd__a21oi_1
X_1386_ net148 net109 net42 VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.data_we\[50\]
+ sky130_fd_sc_hd__and3_2
X_2007_ dig_ctrl_inst.latch_mem_inst.RAM\[57\]\[7\] _0154_ _0160_ dig_ctrl_inst.latch_mem_inst.RAM\[63\]\[7\]
+ VGND VGND VDPWR VDPWR _0712_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_33_362 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[13\].gen_latches\[7\].p_latch net183 dig_ctrl_inst.latch_mem_inst.gclk\[13\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[13\]\[7\] sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[7\].gen_latches\[0\].p_latch net247 dig_ctrl_inst.latch_mem_inst.gclk\[7\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[7\]\[0\] sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_56_498 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_253 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
XFILLER_0_51_234 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[29\].gen_latches\[1\].p_latch net238 dig_ctrl_inst.latch_mem_inst.gclk\[29\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[29\]\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_47_69 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_1240_ net266 dig_ctrl_inst.cpu_inst.r2\[1\] VGND VGND VDPWR VDPWR _1088_ sky130_fd_sc_hd__and2b_1
X_1171_ net258 net254 VGND VGND VDPWR VDPWR _1019_ sky130_fd_sc_hd__or2_4
XFILLER_0_2_27 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XANTENNA_16 ui_in[1] VGND VGND VDPWR VDPWR sky130_fd_sc_hd__diode_2
XANTENNA_27 _1135_ VGND VGND VDPWR VDPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_343 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_125 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_50 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
X_2487_ clknet_leaf_3_clk net333 net173 VGND VGND VDPWR VDPWR dig_ctrl_inst.spi_receiver_inst.spi_sclk_sync
+ sky130_fd_sc_hd__dfrtp_1
X_1507_ _0173_ _0221_ _0216_ dig_ctrl_inst.cpu_inst.ip\[4\] VGND VGND VDPWR VDPWR
+ _0222_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_49_3 VDPWR VGND VDPWR VGND sky130_ef_sc_hd__decap_12
X_1438_ net266 net264 _1020_ _0175_ VGND VGND VDPWR VDPWR _0176_ sky130_fd_sc_hd__nand4_4
X_1369_ net117 net91 net56 VGND VGND VDPWR VDPWR _0141_ sky130_fd_sc_hd__and3_2
XFILLER_0_77_197 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_175 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_337 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_275 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XFILLER_0_68_153 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
Xinput14 uio_in[4] VGND VGND VDPWR VDPWR net14 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_68_197 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_175 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
X_2341_ dig_ctrl_inst.cpu_inst.port_o\[5\] net356 _0986_ VGND VGND VDPWR VDPWR _0092_
+ sky130_fd_sc_hd__mux2_1
X_2410_ clknet_leaf_6_clk _0018_ net145 VGND VGND VDPWR VDPWR dig_ctrl_inst.cpu_inst.port_o\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_58_57 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
X_1154_ dig_ctrl_inst.spi_addr\[2\] VGND VGND VDPWR VDPWR _1003_ sky130_fd_sc_hd__inv_2
X_1223_ net262 dig_ctrl_inst.cpu_inst.r1\[0\] VGND VGND VDPWR VDPWR _1071_ sky130_fd_sc_hd__and2b_1
X_2272_ _0234_ _0785_ _0787_ _0236_ _0957_ VGND VGND VDPWR VDPWR _0958_ sky130_fd_sc_hd__o221ai_1
XFILLER_0_59_164 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
XFILLER_0_59_120 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_337 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[32\].clock_buffer dig_ctrl_inst.latch_mem_inst.gen_gclk\[32\]._gclk
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.gclk\[32\] sky130_fd_sc_hd__clkbuf_4
X_1987_ dig_ctrl_inst.latch_mem_inst.RAM\[35\]\[7\] net131 net102 net51 VGND VGND
+ VDPWR VDPWR _0692_ sky130_fd_sc_hd__and4_1
XFILLER_0_2_194 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_66_560 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout180 dig_ctrl_inst.latch_mem_inst.rst_ni VGND VGND VDPWR VDPWR net180 sky130_fd_sc_hd__clkbuf_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[62\].gen_latches\[1\].p_latch net238 dig_ctrl_inst.latch_mem_inst.gclk\[62\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[62\]\[1\] sky130_fd_sc_hd__dlxtp_1
Xfanout191 net193 VGND VGND VDPWR VDPWR net191 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_72_596 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_25 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_337 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
X_1910_ dig_ctrl_inst.latch_mem_inst.RAM\[34\]\[5\] net109 net52 VGND VGND VDPWR VDPWR
+ _0617_ sky130_fd_sc_hd__and3_2
X_1841_ dig_ctrl_inst.latch_mem_inst.RAM\[4\]\[4\] net123 net97 VGND VGND VDPWR VDPWR
+ _0549_ sky130_fd_sc_hd__and3_2
X_1772_ dig_ctrl_inst.latch_mem_inst.RAM\[21\]\[3\] _0124_ _0478_ _0479_ _0480_ VGND
+ VGND VDPWR VDPWR _0481_ sky130_fd_sc_hd__a2111o_1
X_2324_ _0984_ net355 _0978_ VGND VGND VDPWR VDPWR _0077_ sky130_fd_sc_hd__mux2_1
XFILLER_0_12_248 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_292 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_8
X_1206_ _1018_ _1050_ _1051_ _1052_ _1053_ VGND VGND VDPWR VDPWR _1054_ sky130_fd_sc_hd__o41a_4
X_2186_ _0748_ _0869_ _0875_ _0863_ VGND VGND VDPWR VDPWR _0876_ sky130_fd_sc_hd__o211a_1
X_2255_ _0233_ _0783_ _0936_ _0941_ VGND VGND VDPWR VDPWR _0942_ sky130_fd_sc_hd__a211oi_1
XTAP_TAPCELL_ROW_63_541 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_292 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_101 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_3_185 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_9_Left_87 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_77_633 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2040_ dig_ctrl_inst.cpu_inst.data\[2\] _0449_ _0741_ VGND VGND VDPWR VDPWR _0036_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_60_522 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[63\].clock_gate clknet_leaf_18_clk dig_ctrl_inst.latch_mem_inst.data_we\[63\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.gen_gclk\[63\]._gclk sky130_fd_sc_hd__dlclkp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[55\].gen_latches\[0\].p_latch net242 dig_ctrl_inst.latch_mem_inst.gclk\[55\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[55\]\[0\] sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_17_265 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1755_ _0460_ _0461_ _0462_ _0463_ VGND VGND VDPWR VDPWR _0464_ sky130_fd_sc_hd__or4_2
X_1824_ dig_ctrl_inst.latch_mem_inst.RAM\[37\]\[4\] net117 net100 net54 VGND VGND
+ VDPWR VDPWR _0532_ sky130_fd_sc_hd__and4_1
XFILLER_0_20_61 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
X_1686_ _0287_ _0386_ _0391_ _0396_ VGND VGND VDPWR VDPWR _0397_ sky130_fd_sc_hd__or4_1
X_2238_ dig_ctrl_inst.cpu_inst.r0\[5\] _0758_ _0925_ VGND VGND VDPWR VDPWR _0050_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_29_81 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_2307_ net384 _0975_ _0976_ VGND VGND VDPWR VDPWR _0068_ sky130_fd_sc_hd__mux2_1
XFILLER_0_45_91 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_2169_ _0761_ _0762_ net157 VGND VGND VDPWR VDPWR _0859_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_0_166 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[43\].gen_latches\[7\].p_latch net186 dig_ctrl_inst.latch_mem_inst.gclk\[43\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[43\]\[7\] sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_8_211 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[32\].gen_latches\[5\].p_latch net201 dig_ctrl_inst.latch_mem_inst.gclk\[32\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[32\]\[5\] sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_14_246 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_181 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[21\].gen_latches\[3\].p_latch net215 dig_ctrl_inst.latch_mem_inst.gclk\[21\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[21\]\[3\] sky130_fd_sc_hd__dlxtp_1
X_1540_ _0248_ _0252_ VGND VGND VDPWR VDPWR _0253_ sky130_fd_sc_hd__nand2_1
XFILLER_0_1_215 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_8
X_1471_ dig_ctrl_inst.cpu_inst.r0\[0\] dig_ctrl_inst.cpu_inst.port_o\[0\] _0176_ VGND
+ VGND VDPWR VDPWR _0011_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_49 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_6
Xdig_ctrl_inst.latch_mem_inst.gen_words\[59\].gen_latches\[1\].p_latch net237 dig_ctrl_inst.latch_mem_inst.gclk\[59\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[59\]\[1\] sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_59_Left_137 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
X_2023_ _0710_ _0711_ _0725_ _0727_ VGND VGND VDPWR VDPWR _0728_ sky130_fd_sc_hd__or4_1
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[25\].clock_buffer dig_ctrl_inst.latch_mem_inst.gen_gclk\[25\]._gclk
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.gclk\[25\] sky130_fd_sc_hd__clkbuf_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[10\].gen_latches\[1\].p_latch net235 dig_ctrl_inst.latch_mem_inst.gclk\[10\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[10\]\[1\] sky130_fd_sc_hd__dlxtp_1
X_1807_ dig_ctrl_inst.latch_mem_inst.RAM\[22\]\[4\] net95 net68 VGND VGND VDPWR VDPWR
+ _0515_ sky130_fd_sc_hd__and3_2
XFILLER_0_9_337 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_148 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_68_Left_146 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
X_1738_ _0287_ _0439_ _0442_ _0447_ VGND VGND VDPWR VDPWR _0448_ sky130_fd_sc_hd__or4_4
XFILLER_0_0_281 VDPWR VGND VDPWR VGND sky130_ef_sc_hd__decap_12
X_1669_ dig_ctrl_inst.latch_mem_inst.RAM\[53\]\[1\] _0151_ _0339_ _0340_ _0344_ VGND
+ VGND VDPWR VDPWR _0380_ sky130_fd_sc_hd__a2111o_1
XPHY_EDGE_ROW_77_Left_155 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[3\].gen_latches\[3\].p_latch net220 dig_ctrl_inst.latch_mem_inst.gclk\[3\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[3\]\[3\] sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_36_382 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_232 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[36\].gen_latches\[6\].p_latch net195 dig_ctrl_inst.latch_mem_inst.gclk\[36\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[36\]\[6\] sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_input_latches\[4\].n_latch dig_ctrl_inst.data_out\[4\]
+ clknet_leaf_8_clk VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.wdata\[4\]
+ sky130_fd_sc_hd__dlxtn_2
XFILLER_0_14_129 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[25\].gen_latches\[4\].p_latch net208 dig_ctrl_inst.latch_mem_inst.gclk\[25\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[25\]\[4\] sky130_fd_sc_hd__dlxtp_1
X_1454_ dig_ctrl_inst.spi_addr\[0\] _0186_ VGND VGND VDPWR VDPWR _0187_ sky130_fd_sc_hd__nor2_1
X_1523_ _0234_ _0235_ VGND VGND VDPWR VDPWR _0236_ sky130_fd_sc_hd__or2_1
X_1385_ net156 _0148_ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.data_we\[49\]
+ sky130_fd_sc_hd__and2_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[14\].gen_latches\[2\].p_latch net228 dig_ctrl_inst.latch_mem_inst.gclk\[14\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[14\]\[2\] sky130_fd_sc_hd__dlxtp_1
X_2006_ dig_ctrl_inst.latch_mem_inst.RAM\[10\]\[7\] net123 net294 _0700_ _0709_ VGND
+ VGND VDPWR VDPWR _0711_ sky130_fd_sc_hd__a311o_1
XTAP_TAPCELL_ROW_33_363 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[7\].gen_latches\[4\].p_latch net212 dig_ctrl_inst.latch_mem_inst.gclk\[7\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[7\]\[4\] sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_56_499 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_287 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_15 VDPWR VGND VDPWR VGND sky130_ef_sc_hd__decap_12
X_1170_ net258 net254 VGND VGND VDPWR VDPWR _1018_ sky130_fd_sc_hd__nor2_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[29\].gen_latches\[5\].p_latch net204 dig_ctrl_inst.latch_mem_inst.gclk\[29\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[29\]\[5\] sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_47_444 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_28 dig_ctrl_inst.cpu_inst.port_o\[5\] VGND VGND VDPWR VDPWR sky130_fd_sc_hd__diode_2
XANTENNA_17 ui_in[3] VGND VGND VDPWR VDPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_344 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2486_ clknet_leaf_3_clk net13 net173 VGND VGND VDPWR VDPWR dig_ctrl_inst.spi_receiver_inst.synchronizer_spi_sclk.pipe\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_1437_ dig_ctrl_inst.cpu_inst.skip _0174_ VGND VGND VDPWR VDPWR _0175_ sky130_fd_sc_hd__nor2_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[18\].gen_latches\[3\].p_latch net219 dig_ctrl_inst.latch_mem_inst.gclk\[18\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[18\]\[3\] sky130_fd_sc_hd__dlxtp_1
X_1506_ net159 dig_ctrl_inst.cpu_inst.data\[4\] _0198_ VGND VGND VDPWR VDPWR _0221_
+ sky130_fd_sc_hd__mux2_1
X_1299_ net155 _1139_ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.data_we\[7\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_37_70 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
X_1368_ net149 net86 net53 VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.data_we\[40\]
+ sky130_fd_sc_hd__and3_2
XFILLER_0_18_287 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_290 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_181 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_69_580 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_18 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_6
Xinput15 uio_in[5] VGND VGND VDPWR VDPWR net15 sky130_fd_sc_hd__buf_1
X_2340_ dig_ctrl_inst.cpu_inst.port_o\[4\] net348 _0986_ VGND VGND VDPWR VDPWR _0091_
+ sky130_fd_sc_hd__mux2_1
X_2271_ _0786_ _0791_ _0172_ VGND VGND VDPWR VDPWR _0957_ sky130_fd_sc_hd__mux2_1
XFILLER_0_74_79 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_1153_ net251 VGND VGND VDPWR VDPWR _1002_ sky130_fd_sc_hd__inv_2
X_1222_ net265 dig_ctrl_inst.cpu_inst.r2\[0\] VGND VGND VDPWR VDPWR _1070_ sky130_fd_sc_hd__and2b_1
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[18\].clock_buffer dig_ctrl_inst.latch_mem_inst.gen_gclk\[18\]._gclk
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.gclk\[18\] sky130_fd_sc_hd__clkbuf_4
X_1986_ dig_ctrl_inst.latch_mem_inst.RAM\[60\]\[7\] net78 net48 VGND VGND VDPWR VDPWR
+ _0691_ sky130_fd_sc_hd__and3_2
XFILLER_0_47_327 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_9_clk clknet_1_1__leaf_clk VGND VGND VDPWR VDPWR clknet_leaf_9_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_15_235 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_246 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_279 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_2469_ clknet_leaf_10_clk _0075_ net142 VGND VGND VDPWR VDPWR dig_ctrl_inst.cpu_inst.r3\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_66_561 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_113 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_305 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_341 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
Xfanout181 _1021_ VGND VGND VDPWR VDPWR net181 sky130_fd_sc_hd__buf_6
XFILLER_0_44_27 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
Xfanout170 net171 VGND VGND VDPWR VDPWR net170 sky130_fd_sc_hd__buf_2
Xfanout192 net193 VGND VGND VDPWR VDPWR net192 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_TAPCELL_ROW_72_597 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[62\].gen_latches\[5\].p_latch net205 dig_ctrl_inst.latch_mem_inst.gclk\[62\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[62\]\[5\] sky130_fd_sc_hd__dlxtp_1
X_1840_ dig_ctrl_inst.latch_mem_inst.RAM\[18\]\[4\] net111 net68 VGND VGND VDPWR VDPWR
+ _0548_ sky130_fd_sc_hd__and3_2
XFILLER_0_69_57 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_341 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_31_Left_109 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
X_1771_ dig_ctrl_inst.latch_mem_inst.RAM\[31\]\[3\] net103 net80 net62 VGND VGND VDPWR
+ VDPWR _0480_ sky130_fd_sc_hd__and4_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[51\].gen_latches\[3\].p_latch net222 dig_ctrl_inst.latch_mem_inst.gclk\[51\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[51\]\[3\] sky130_fd_sc_hd__dlxtp_1
X_2323_ dig_ctrl_inst.spi_receiver_inst.spi_cnt\[2\] _0979_ _0981_ _0983_ VGND VGND
+ VDPWR VDPWR _0984_ sky130_fd_sc_hd__o22a_1
X_2254_ _0937_ _0938_ _0940_ VGND VGND VDPWR VDPWR _0941_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_63_542 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1205_ net260 net256 dig_ctrl_inst.cpu_inst.r0\[2\] VGND VGND VDPWR VDPWR _1053_
+ sky130_fd_sc_hd__or3_1
XPHY_EDGE_ROW_40_Left_118 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
X_2185_ _0870_ _0871_ _0874_ VGND VGND VDPWR VDPWR _0875_ sky130_fd_sc_hd__and3_2
XFILLER_0_18_83 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_341 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
Xclone18 _1021_ VGND VGND VDPWR VDPWR net300 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_7_232 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_254 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_287 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
X_1969_ dig_ctrl_inst.latch_mem_inst.RAM\[33\]\[6\] _0135_ _0632_ _0633_ _0639_ VGND
+ VGND VDPWR VDPWR _0675_ sky130_fd_sc_hd__a2111o_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[40\].gen_latches\[1\].p_latch net234 dig_ctrl_inst.latch_mem_inst.gclk\[40\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[40\]\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_11_260 VDPWR VGND VDPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_634 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_523 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_135 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_113 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_1823_ dig_ctrl_inst.latch_mem_inst.RAM\[42\]\[4\] net84 net54 VGND VGND VDPWR VDPWR
+ _0531_ sky130_fd_sc_hd__and3_2
XTAP_TAPCELL_ROW_17_266 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[55\].gen_latches\[4\].p_latch net208 dig_ctrl_inst.latch_mem_inst.gclk\[55\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[55\]\[4\] sky130_fd_sc_hd__dlxtp_1
X_1754_ dig_ctrl_inst.latch_mem_inst.RAM\[12\]\[3\] _1148_ _0129_ dig_ctrl_inst.latch_mem_inst.RAM\[26\]\[3\]
+ VGND VGND VDPWR VDPWR _0463_ sky130_fd_sc_hd__a22o_1
Xmax_cap134 _1094_ VGND VGND VDPWR VDPWR net134 sky130_fd_sc_hd__buf_4
XFILLER_0_4_235 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_1685_ _0392_ _0393_ _0394_ _0395_ VGND VGND VDPWR VDPWR _0396_ sky130_fd_sc_hd__or4_1
X_2237_ _0920_ _0924_ VGND VGND VDPWR VDPWR _0925_ sky130_fd_sc_hd__nand2b_1
X_2306_ net363 _0974_ _0976_ VGND VGND VDPWR VDPWR _0067_ sky130_fd_sc_hd__mux2_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[44\].gen_latches\[2\].p_latch net226 dig_ctrl_inst.latch_mem_inst.gclk\[44\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[44\]\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_24_3 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
X_2168_ dig_ctrl_inst.cpu_inst.r0\[3\] net41 VGND VGND VDPWR VDPWR _0858_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_0_167 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_156 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2099_ _1016_ _0745_ VGND VGND VDPWR VDPWR _0792_ sky130_fd_sc_hd__nor2_1
XFILLER_0_43_182 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[33\].gen_latches\[0\].p_latch net240 dig_ctrl_inst.latch_mem_inst.gclk\[33\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[33\]\[0\] sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_17_Right_17 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_26_Right_26 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_8_212 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_18 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_35_Right_35 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_138 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_14_247 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1470_ dig_ctrl_inst.spi_addr\[5\] _0196_ _0197_ VGND VGND VDPWR VDPWR _0010_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_1_238 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_6
Xdig_ctrl_inst.latch_mem_inst.gen_words\[21\].gen_latches\[7\].p_latch net183 dig_ctrl_inst.latch_mem_inst.gclk\[21\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[21\]\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_66_58 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_44_Right_44 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_39 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[10\].gen_latches\[5\].p_latch net204 dig_ctrl_inst.latch_mem_inst.gclk\[10\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[10\]\[5\] sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[59\].gen_latches\[5\].p_latch net204 dig_ctrl_inst.latch_mem_inst.gclk\[59\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[59\]\[5\] sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_53_Right_53 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
X_2022_ _0712_ _0726_ VGND VGND VDPWR VDPWR _0727_ sky130_fd_sc_hd__or2_1
XFILLER_0_9_327 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_1806_ dig_ctrl_inst.latch_mem_inst.RAM\[20\]\[4\] net97 net68 VGND VGND VDPWR VDPWR
+ _0514_ sky130_fd_sc_hd__and3_2
XFILLER_0_31_83 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_193 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_62_Right_62 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
X_1737_ _0443_ _0444_ _0445_ _0446_ VGND VGND VDPWR VDPWR _0447_ sky130_fd_sc_hd__or4_1
X_1599_ dig_ctrl_inst.latch_mem_inst.RAM\[56\]\[0\] net87 net45 _0146_ dig_ctrl_inst.latch_mem_inst.RAM\[47\]\[0\]
+ VGND VGND VDPWR VDPWR _0311_ sky130_fd_sc_hd__a32o_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[48\].gen_latches\[3\].p_latch net215 dig_ctrl_inst.latch_mem_inst.gclk\[48\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[48\]\[3\] sky130_fd_sc_hd__dlxtp_1
X_1668_ dig_ctrl_inst.latch_mem_inst.RAM\[33\]\[1\] _0135_ _0352_ _0369_ _0372_ VGND
+ VGND VDPWR VDPWR _0379_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_0_293 VDPWR VGND VDPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_71_Right_71 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[3\].gen_latches\[7\].p_latch net187 dig_ctrl_inst.latch_mem_inst.gclk\[3\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[3\]\[7\] sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_36_383 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_228 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[37\].gen_latches\[1\].p_latch net234 dig_ctrl_inst.latch_mem_inst.gclk\[37\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[37\]\[1\] sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_12_Left_90 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_244 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_46 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_1453_ net251 dig_ctrl_inst.mode_d dig_ctrl_inst.spi_receiver_inst.stb_o VGND VGND
+ VDPWR VDPWR _0186_ sky130_fd_sc_hd__and3_2
X_1522_ _0172_ _0233_ VGND VGND VDPWR VDPWR _0235_ sky130_fd_sc_hd__and2_1
XFILLER_0_22_141 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
X_1384_ net132 net118 net50 VGND VGND VDPWR VDPWR _0148_ sky130_fd_sc_hd__and3_2
X_2005_ dig_ctrl_inst.latch_mem_inst.RAM\[44\]\[7\] _0144_ _0159_ dig_ctrl_inst.latch_mem_inst.RAM\[62\]\[7\]
+ _0701_ VGND VGND VDPWR VDPWR _0710_ sky130_fd_sc_hd__a221o_1
XFILLER_0_26_50 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[14\].gen_latches\[6\].p_latch net192 dig_ctrl_inst.latch_mem_inst.gclk\[14\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[14\]\[6\] sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_33_364 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_341 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_185 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_277 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_211 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_47_445 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_29 VDPWR VGND VDPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_18 ui_in[7] VGND VGND VDPWR VDPWR sky130_fd_sc_hd__diode_2
XFILLER_0_59_314 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
XANTENNA_29 dig_ctrl_inst.latch_mem_inst.gclk\[19\] VGND VGND VDPWR VDPWR sky130_fd_sc_hd__diode_2
XFILLER_0_42_247 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_30_345 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2485_ clknet_leaf_3_clk net337 net176 VGND VGND VDPWR VDPWR dig_ctrl_inst.spi_receiver_inst.spi_cs_sync
+ sky130_fd_sc_hd__dfrtp_1
X_1436_ net248 dig_ctrl_inst.cpu_inst.cpu_state\[1\] _0999_ VGND VGND VDPWR VDPWR
+ _0174_ sky130_fd_sc_hd__nand3_2
X_1505_ _0204_ _0219_ VGND VGND VDPWR VDPWR _0220_ sky130_fd_sc_hd__or2_1
XFILLER_0_10_166 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
X_1367_ net86 net53 VGND VGND VDPWR VDPWR _0140_ sky130_fd_sc_hd__and2_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[18\].gen_latches\[7\].p_latch net186 dig_ctrl_inst.latch_mem_inst.gclk\[18\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[18\]\[7\] sky130_fd_sc_hd__dlxtp_1
X_1298_ net126 net106 net101 VGND VGND VDPWR VDPWR _1139_ sky130_fd_sc_hd__and3_2
XFILLER_0_33_236 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_225 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_299 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_69_581 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_166 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_44_426 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[57\].clock_buffer dig_ctrl_inst.latch_mem_inst.gen_gclk\[57\]._gclk
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.gclk\[57\] sky130_fd_sc_hd__clkbuf_4
X_2270_ _0233_ _0933_ VGND VGND VDPWR VDPWR _0956_ sky130_fd_sc_hd__xnor2_1
X_1221_ net265 net262 dig_ctrl_inst.cpu_inst.r3\[0\] VGND VGND VDPWR VDPWR _1069_
+ sky130_fd_sc_hd__and3_2
XFILLER_0_59_133 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_1152_ dig_ctrl_inst.cpu_inst.ip\[0\] VGND VGND VDPWR VDPWR _1001_ sky130_fd_sc_hd__inv_2
X_1985_ dig_ctrl_inst.latch_mem_inst.RAM\[29\]\[7\] net118 net82 net69 VGND VGND VDPWR
+ VDPWR _0690_ sky130_fd_sc_hd__and4_1
XFILLER_0_23_84 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_174 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
X_2399_ clknet_leaf_3_clk _0008_ net172 VGND VGND VDPWR VDPWR dig_ctrl_inst.spi_addr\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_1419_ net249 dig_ctrl_inst.spi_data_o\[4\] _1118_ _0162_ VGND VGND VDPWR VDPWR dig_ctrl_inst.data_out\[4\]
+ sky130_fd_sc_hd__a22o_1
X_2468_ clknet_leaf_7_clk _0074_ net144 VGND VGND VDPWR VDPWR dig_ctrl_inst.cpu_inst.r3\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_66_562 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire40 _0459_ VGND VGND VDPWR VDPWR net40 sky130_fd_sc_hd__clkbuf_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[63\].gen_latches\[0\].p_latch net242 dig_ctrl_inst.latch_mem_inst.gclk\[63\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[63\]\[0\] sky130_fd_sc_hd__dlxtp_1
Xfanout193 net194 VGND VGND VDPWR VDPWR net193 sky130_fd_sc_hd__clkbuf_2
Xfanout171 _1036_ VGND VGND VDPWR VDPWR net171 sky130_fd_sc_hd__clkbuf_2
Xfanout160 _1110_ VGND VGND VDPWR VDPWR net160 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_72_598 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_169 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_1770_ dig_ctrl_inst.latch_mem_inst.RAM\[50\]\[3\] net110 net44 VGND VGND VDPWR VDPWR
+ _0479_ sky130_fd_sc_hd__and3_2
XFILLER_0_69_36 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_2322_ dig_ctrl_inst.spi_receiver_inst.spi_cnt\[1\] _0982_ dig_ctrl_inst.spi_receiver_inst.spi_cnt\[2\]
+ VGND VGND VDPWR VDPWR _0983_ sky130_fd_sc_hd__a21bo_1
X_1204_ net256 dig_ctrl_inst.cpu_inst.r1\[2\] VGND VGND VDPWR VDPWR _1052_ sky130_fd_sc_hd__and2b_1
X_2184_ _0749_ _0869_ _0873_ VGND VGND VDPWR VDPWR _0874_ sky130_fd_sc_hd__a21oi_1
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[14\].clock_gate clknet_leaf_17_clk dig_ctrl_inst.latch_mem_inst.data_we\[14\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.gen_gclk\[14\]._gclk sky130_fd_sc_hd__dlclkp_1
X_2253_ _0230_ _0787_ _0939_ VGND VGND VDPWR VDPWR _0940_ sky130_fd_sc_hd__o21ai_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[51\].gen_latches\[7\].p_latch net183 dig_ctrl_inst.latch_mem_inst.gclk\[51\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[51\]\[7\] sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_63_543 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1968_ _0673_ _0665_ _0672_ _0664_ VGND VGND VDPWR VDPWR _0674_ sky130_fd_sc_hd__or4_4
XFILLER_0_50_71 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_8
Xdig_ctrl_inst.latch_mem_inst.gen_words\[40\].gen_latches\[5\].p_latch net202 dig_ctrl_inst.latch_mem_inst.gclk\[40\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[40\]\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_7_222 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_266 VDPWR VGND VDPWR VGND sky130_ef_sc_hd__decap_12
X_1899_ dig_ctrl_inst.latch_mem_inst.RAM\[32\]\[5\] net128 net55 VGND VGND VDPWR VDPWR
+ _0606_ sky130_fd_sc_hd__and3_2
XFILLER_0_11_272 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_161 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_77_635 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_624 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_267 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1753_ dig_ctrl_inst.latch_mem_inst.RAM\[15\]\[3\] _0117_ _0142_ dig_ctrl_inst.latch_mem_inst.RAM\[42\]\[3\]
+ VGND VGND VDPWR VDPWR _0462_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_60_524 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1822_ dig_ctrl_inst.latch_mem_inst.RAM\[63\]\[4\] net104 net81 net45 VGND VGND VDPWR
+ VDPWR _0530_ sky130_fd_sc_hd__and4_1
XFILLER_0_52_194 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
X_1684_ dig_ctrl_inst.latch_mem_inst.RAM\[41\]\[1\] _0141_ _0347_ _0351_ _0362_ VGND
+ VGND VDPWR VDPWR _0395_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_20_85 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_96 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
X_2236_ _0754_ _0922_ _0923_ _0756_ net41 VGND VGND VDPWR VDPWR _0924_ sky130_fd_sc_hd__o221a_1
X_2167_ dig_ctrl_inst.cpu_inst.r0\[2\] _0857_ _0758_ VGND VGND VDPWR VDPWR _0047_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_45_71 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
X_2305_ net366 _0973_ _0976_ VGND VGND VDPWR VDPWR _0066_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_3 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[44\].gen_latches\[6\].p_latch net197 dig_ctrl_inst.latch_mem_inst.gclk\[44\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[44\]\[6\] sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[0\].gen_latches\[1\].p_latch net239 dig_ctrl_inst.latch_mem_inst.gclk\[0\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[0\]\[1\] sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_0_157 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2098_ _1016_ _0744_ VGND VGND VDPWR VDPWR _0791_ sky130_fd_sc_hd__or2_1
XFILLER_0_16_331 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_8
Xdig_ctrl_inst.latch_mem_inst.gen_words\[33\].gen_latches\[4\].p_latch net210 dig_ctrl_inst.latch_mem_inst.gclk\[33\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[33\]\[4\] sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_8_213 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[22\].gen_latches\[2\].p_latch net226 dig_ctrl_inst.latch_mem_inst.gclk\[22\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[22\]\[2\] sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_14_248 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_15 VDPWR VGND VDPWR VGND sky130_ef_sc_hd__decap_12
Xdig_ctrl_inst.latch_mem_inst.gen_words\[11\].gen_latches\[0\].p_latch net243 dig_ctrl_inst.latch_mem_inst.gclk\[11\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[11\]\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_34_194 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
X_2021_ dig_ctrl_inst.latch_mem_inst.RAM\[28\]\[7\] net77 net65 _0127_ dig_ctrl_inst.latch_mem_inst.RAM\[24\]\[7\]
+ VGND VGND VDPWR VDPWR _0726_ sky130_fd_sc_hd__a32o_1
X_1805_ dig_ctrl_inst.latch_mem_inst.RAM\[32\]\[4\] _0134_ _0148_ dig_ctrl_inst.latch_mem_inst.RAM\[49\]\[4\]
+ VGND VGND VDPWR VDPWR _0513_ sky130_fd_sc_hd__a22o_1
X_1736_ dig_ctrl_inst.latch_mem_inst.RAM\[49\]\[2\] _0148_ _0400_ _0411_ _0413_ VGND
+ VGND VDPWR VDPWR _0446_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_40_153 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
X_1667_ dig_ctrl_inst.latch_mem_inst.RAM\[1\]\[1\] _1130_ _1148_ dig_ctrl_inst.latch_mem_inst.RAM\[12\]\[1\]
+ VGND VGND VDPWR VDPWR _0378_ sky130_fd_sc_hd__a22o_1
X_1598_ dig_ctrl_inst.latch_mem_inst.RAM\[22\]\[0\] _0125_ _0154_ dig_ctrl_inst.latch_mem_inst.RAM\[57\]\[0\]
+ VGND VGND VDPWR VDPWR _0310_ sky130_fd_sc_hd__a22o_1
XFILLER_0_40_186 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_164 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_6
Xdig_ctrl_inst.latch_mem_inst.gen_words\[4\].gen_latches\[2\].p_latch net229 dig_ctrl_inst.latch_mem_inst.gclk\[4\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[4\]\[2\] sky130_fd_sc_hd__dlxtp_1
X_2219_ _0244_ _0906_ VGND VGND VDPWR VDPWR _0907_ sky130_fd_sc_hd__xnor2_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[48\].gen_latches\[7\].p_latch net183 dig_ctrl_inst.latch_mem_inst.gclk\[48\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[48\]\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_48_242 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[37\].gen_latches\[5\].p_latch net203 dig_ctrl_inst.latch_mem_inst.gclk\[37\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[37\]\[5\] sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_11_229 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_150 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_142 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_3 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_8
Xdig_ctrl_inst.latch_mem_inst.gen_words\[26\].gen_latches\[3\].p_latch net222 dig_ctrl_inst.latch_mem_inst.gclk\[26\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[26\]\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_39_275 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_309 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[15\].gen_latches\[1\].p_latch net235 dig_ctrl_inst.latch_mem_inst.gclk\[15\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[15\]\[1\] sky130_fd_sc_hd__dlxtp_1
X_1452_ _1096_ _0184_ VGND VGND VDPWR VDPWR _0185_ sky130_fd_sc_hd__nand2_1
X_1383_ net128 net150 net44 VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.data_we\[48\]
+ sky130_fd_sc_hd__and3_2
XFILLER_0_10_337 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
X_1521_ _0172_ _0233_ VGND VGND VDPWR VDPWR _0234_ sky130_fd_sc_hd__nor2_1
XFILLER_0_77_315 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_2004_ dig_ctrl_inst.latch_mem_inst.RAM\[1\]\[7\] _1130_ _0138_ dig_ctrl_inst.latch_mem_inst.RAM\[37\]\[7\]
+ VGND VGND VDPWR VDPWR _0709_ sky130_fd_sc_hd__a22o_1
XFILLER_0_42_83 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_33_365 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_169 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[8\].gen_latches\[3\].p_latch net217 dig_ctrl_inst.latch_mem_inst.gclk\[8\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[8\]\[3\] sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[21\].clock_buffer dig_ctrl_inst.latch_mem_inst.gen_gclk\[21\]._gclk
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.gclk\[21\] sky130_fd_sc_hd__clkbuf_4
X_1719_ dig_ctrl_inst.latch_mem_inst.RAM\[16\]\[2\] _0119_ _0146_ dig_ctrl_inst.latch_mem_inst.RAM\[47\]\[2\]
+ _0428_ VGND VGND VDPWR VDPWR _0429_ sky130_fd_sc_hd__a221o_1
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[7\].clock_buffer dig_ctrl_inst.latch_mem_inst.gen_gclk\[7\]._gclk
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.gclk\[7\] sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_24_310 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[19\].clock_gate clknet_leaf_0_clk dig_ctrl_inst.latch_mem_inst.data_we\[19\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.gen_gclk\[19\]._gclk sky130_fd_sc_hd__dlclkp_1
XFILLER_0_59_337 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_47_446 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_19 uio_in[0] VGND VGND VDPWR VDPWR sky130_fd_sc_hd__diode_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[19\].gen_latches\[2\].p_latch net229 dig_ctrl_inst.latch_mem_inst.gclk\[19\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[19\]\[2\] sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_30_346 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_245 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_223 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_201 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_20 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
X_1504_ dig_ctrl_inst.cpu_inst.ip\[4\] _0215_ _0173_ VGND VGND VDPWR VDPWR _0219_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_2_312 VDPWR VGND VDPWR VGND sky130_ef_sc_hd__decap_12
X_2484_ clknet_leaf_3_clk net11 net173 VGND VGND VDPWR VDPWR dig_ctrl_inst.spi_receiver_inst.synchronizer_spi_cs.pipe\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_1366_ net156 _0139_ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.data_we\[39\]
+ sky130_fd_sc_hd__and2_1
X_1435_ net248 dig_ctrl_inst.cpu_inst.cpu_state\[1\] _0999_ VGND VGND VDPWR VDPWR
+ _0173_ sky130_fd_sc_hd__and3_2
X_1297_ net148 net120 net93 VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.data_we\[6\]
+ sky130_fd_sc_hd__and3_2
XFILLER_0_5_161 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[21\].clock_gate clknet_leaf_15_clk dig_ctrl_inst.latch_mem_inst.data_we\[21\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.gen_gclk\[21\]._gclk sky130_fd_sc_hd__dlclkp_1
XTAP_TAPCELL_ROW_44_427 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_19 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
X_1151_ net254 VGND VGND VDPWR VDPWR _1000_ sky130_fd_sc_hd__inv_2
X_1220_ net157 VGND VGND VDPWR VDPWR _1068_ sky130_fd_sc_hd__inv_2
X_1984_ dig_ctrl_inst.latch_mem_inst.RAM\[12\]\[7\] net122 net76 VGND VGND VDPWR VDPWR
+ _0689_ sky130_fd_sc_hd__and3_2
X_2467_ clknet_leaf_7_clk _0073_ net143 VGND VGND VDPWR VDPWR dig_ctrl_inst.cpu_inst.r3\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_197 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
X_1349_ net153 net73 net70 VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.data_we\[30\]
+ sky130_fd_sc_hd__and3_2
XTAP_TAPCELL_ROW_66_563 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2398_ clknet_leaf_2_clk _0007_ net172 VGND VGND VDPWR VDPWR dig_ctrl_inst.spi_addr\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_1418_ net249 dig_ctrl_inst.spi_data_o\[3\] _1036_ _0162_ VGND VGND VDPWR VDPWR dig_ctrl_inst.data_out\[3\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_47_3 VDPWR VGND VDPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_408 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout172 net176 VGND VGND VDPWR VDPWR net172 sky130_fd_sc_hd__clkbuf_4
Xfanout161 _1090_ VGND VGND VDPWR VDPWR net161 sky130_fd_sc_hd__buf_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[63\].gen_latches\[4\].p_latch net209 dig_ctrl_inst.latch_mem_inst.gclk\[63\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[63\]\[4\] sky130_fd_sc_hd__dlxtp_1
Xfanout150 net151 VGND VGND VDPWR VDPWR net150 sky130_fd_sc_hd__clkbuf_2
Xfanout183 net184 VGND VGND VDPWR VDPWR net183 sky130_fd_sc_hd__clkbuf_2
Xfanout194 net322 VGND VGND VDPWR VDPWR net194 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_72_599 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_17 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_29 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[52\].gen_latches\[2\].p_latch net225 dig_ctrl_inst.latch_mem_inst.gclk\[52\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[52\]\[2\] sky130_fd_sc_hd__dlxtp_1
X_2321_ dig_ctrl_inst.spi_data_i\[1\] dig_ctrl_inst.spi_data_i\[0\] dig_ctrl_inst.spi_receiver_inst.spi_cnt\[0\]
+ VGND VGND VDPWR VDPWR _0982_ sky130_fd_sc_hd__mux2_1
XFILLER_0_69_26 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_251 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_1203_ net260 net256 dig_ctrl_inst.cpu_inst.r3\[2\] VGND VGND VDPWR VDPWR _1051_
+ sky130_fd_sc_hd__and3_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[41\].gen_latches\[0\].p_latch net240 dig_ctrl_inst.latch_mem_inst.gclk\[41\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[41\]\[0\] sky130_fd_sc_hd__dlxtp_1
X_2183_ net159 _0783_ _0790_ net170 _0872_ VGND VGND VDPWR VDPWR _0873_ sky130_fd_sc_hd__a221o_1
X_2252_ _0786_ _0791_ _0167_ VGND VGND VDPWR VDPWR _0939_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_63_544 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_340 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_192 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
X_1967_ _0137_ dig_ctrl_inst.latch_mem_inst.RAM\[35\]\[6\] _0635_ _0642_ _0650_ VGND
+ VGND VDPWR VDPWR _0673_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_7_278 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
X_1898_ dig_ctrl_inst.latch_mem_inst.RAM\[14\]\[5\] net120 net72 VGND VGND VDPWR VDPWR
+ _0605_ sky130_fd_sc_hd__and3_2
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[14\].clock_buffer dig_ctrl_inst.latch_mem_inst.gen_gclk\[14\]._gclk
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.gclk\[14\] sky130_fd_sc_hd__clkbuf_4
X_2519_ net269 VGND VGND VDPWR VDPWR uio_oe[0] sky130_fd_sc_hd__buf_2
XFILLER_0_11_251 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_77_625 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_525 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[56\].gen_latches\[3\].p_latch net218 dig_ctrl_inst.latch_mem_inst.gclk\[56\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[56\]\[3\] sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_17_268 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1752_ dig_ctrl_inst.latch_mem_inst.RAM\[28\]\[3\] net79 net69 _0155_ dig_ctrl_inst.latch_mem_inst.RAM\[58\]\[3\]
+ VGND VGND VDPWR VDPWR _0461_ sky130_fd_sc_hd__a32o_1
Xclkbuf_leaf_10_clk clknet_1_0__leaf_clk VGND VGND VDPWR VDPWR clknet_leaf_10_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_4_215 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
X_1683_ dig_ctrl_inst.latch_mem_inst.RAM\[9\]\[1\] _1143_ _0349_ _0357_ _0361_ VGND
+ VGND VDPWR VDPWR _0394_ sky130_fd_sc_hd__a2111o_1
X_1821_ dig_ctrl_inst.latch_mem_inst.RAM\[40\]\[4\] _0140_ _0153_ dig_ctrl_inst.latch_mem_inst.RAM\[55\]\[4\]
+ _0528_ VGND VGND VDPWR VDPWR _0529_ sky130_fd_sc_hd__a221o_1
Xmax_cap136 _1048_ VGND VGND VDPWR VDPWR net136 sky130_fd_sc_hd__buf_6
X_2304_ net378 _0972_ _0976_ VGND VGND VDPWR VDPWR _0065_ sky130_fd_sc_hd__mux2_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[45\].gen_latches\[1\].p_latch net234 dig_ctrl_inst.latch_mem_inst.gclk\[45\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[45\]\[1\] sky130_fd_sc_hd__dlxtp_1
X_2235_ dig_ctrl_inst.synchronizer_port_i_inst\[5\].out _0802_ _0804_ dig_ctrl_inst.spi_data_o\[5\]
+ VGND VGND VDPWR VDPWR _0923_ sky130_fd_sc_hd__a22oi_1
X_2166_ _0756_ _0855_ _0856_ _0754_ _0854_ VGND VGND VDPWR VDPWR _0857_ sky130_fd_sc_hd__o221ai_1
XTAP_TAPCELL_ROW_0_158 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2097_ _1016_ _0744_ VGND VGND VDPWR VDPWR _0790_ sky130_fd_sc_hd__nor2_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[0\].gen_latches\[5\].p_latch net207 dig_ctrl_inst.latch_mem_inst.gclk\[0\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[0\]\[5\] sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[0\].clock_gate clknet_leaf_9_clk dig_ctrl_inst.latch_mem_inst.data_we\[0\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.gen_gclk\[0\]._gclk sky130_fd_sc_hd__dlclkp_1
XPHY_EDGE_ROW_3_Right_3 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_41 VDPWR VGND VDPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_214 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_74_606 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_1__f_clk clknet_0_clk VGND VGND VDPWR VDPWR clknet_1_1__leaf_clk sky130_fd_sc_hd__clkbuf_16
Xdig_ctrl_inst.latch_mem_inst.gen_words\[22\].gen_latches\[6\].p_latch net197 dig_ctrl_inst.latch_mem_inst.gclk\[22\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[22\]\[6\] sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_14_249 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_324 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_27 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_19 VDPWR VGND VDPWR VGND sky130_ef_sc_hd__decap_12
Xdig_ctrl_inst.latch_mem_inst.gen_words\[11\].gen_latches\[4\].p_latch net214 dig_ctrl_inst.latch_mem_inst.gclk\[11\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[11\]\[4\] sky130_fd_sc_hd__dlxtp_1
X_2020_ dig_ctrl_inst.latch_mem_inst.RAM\[14\]\[7\] _0116_ _0140_ dig_ctrl_inst.latch_mem_inst.RAM\[40\]\[7\]
+ _0713_ VGND VGND VDPWR VDPWR _0725_ sky130_fd_sc_hd__a221o_1
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[26\].clock_gate clknet_leaf_0_clk dig_ctrl_inst.latch_mem_inst.data_we\[26\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.gen_gclk\[26\]._gclk sky130_fd_sc_hd__dlclkp_1
XFILLER_0_57_276 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_28_Left_106 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
X_1735_ dig_ctrl_inst.latch_mem_inst.RAM\[13\]\[2\] _0114_ _0405_ _0414_ _0416_ VGND
+ VGND VDPWR VDPWR _0445_ sky130_fd_sc_hd__a2111o_1
X_1666_ dig_ctrl_inst.latch_mem_inst.RAM\[58\]\[1\] _0155_ _0159_ dig_ctrl_inst.latch_mem_inst.RAM\[62\]\[1\]
+ VGND VGND VDPWR VDPWR _0377_ sky130_fd_sc_hd__a22o_1
X_1804_ dig_ctrl_inst.latch_mem_inst.RAM\[3\]\[4\] _1135_ _0149_ dig_ctrl_inst.latch_mem_inst.RAM\[51\]\[4\]
+ VGND VGND VDPWR VDPWR _0512_ sky130_fd_sc_hd__a22o_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[49\].gen_latches\[2\].p_latch net228 dig_ctrl_inst.latch_mem_inst.gclk\[49\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[49\]\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_40_176 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
X_1597_ dig_ctrl_inst.latch_mem_inst.RAM\[38\]\[0\] net95 net57 _0145_ dig_ctrl_inst.latch_mem_inst.RAM\[45\]\[0\]
+ VGND VGND VDPWR VDPWR _0309_ sky130_fd_sc_hd__a32o_1
XPHY_EDGE_ROW_37_Left_115 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[38\].gen_latches\[0\].p_latch net244 dig_ctrl_inst.latch_mem_inst.gclk\[38\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[38\]\[0\] sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[4\].gen_latches\[6\].p_latch net198 dig_ctrl_inst.latch_mem_inst.gclk\[4\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[4\]\[6\] sky130_fd_sc_hd__dlxtp_1
X_2149_ _0768_ _0780_ VGND VGND VDPWR VDPWR _0840_ sky130_fd_sc_hd__or2_1
X_2218_ _0240_ _0884_ _0238_ VGND VGND VDPWR VDPWR _0906_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_63_279 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_46_Left_124 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_55_Left_133 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[26\].gen_latches\[7\].p_latch net188 dig_ctrl_inst.latch_mem_inst.gclk\[26\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[26\]\[7\] sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_64_Left_142 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_29 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_26 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_73_Left_151 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
X_1520_ net265 net262 dig_ctrl_inst.cpu_inst.r0\[7\] _0231_ _0232_ VGND VGND VDPWR
+ VDPWR _0233_ sky130_fd_sc_hd__o32a_4
X_1451_ _1002_ dig_ctrl_inst.mode_d VGND VGND VDPWR VDPWR _0184_ sky130_fd_sc_hd__or2_1
X_1382_ _1112_ _1127_ VGND VGND VDPWR VDPWR _0147_ sky130_fd_sc_hd__and2_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[15\].gen_latches\[5\].p_latch net199 dig_ctrl_inst.latch_mem_inst.gclk\[15\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[15\]\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_10_327 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
X_2003_ dig_ctrl_inst.latch_mem_inst.RAM\[30\]\[7\] net74 net69 VGND VGND VDPWR VDPWR
+ _0708_ sky130_fd_sc_hd__and3_2
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[60\].clock_buffer dig_ctrl_inst.latch_mem_inst.gen_gclk\[60\]._gclk
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.gclk\[60\] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_5_310 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
XFILLER_0_77_3 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_40 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_8
X_1649_ dig_ctrl_inst.latch_mem_inst.RAM\[37\]\[1\] net115 net99 net52 VGND VGND VDPWR
+ VDPWR _0360_ sky130_fd_sc_hd__and4_1
X_1718_ dig_ctrl_inst.latch_mem_inst.RAM\[2\]\[2\] _1133_ _0152_ dig_ctrl_inst.latch_mem_inst.RAM\[54\]\[2\]
+ VGND VGND VDPWR VDPWR _0428_ sky130_fd_sc_hd__a22o_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[8\].gen_latches\[7\].p_latch net187 dig_ctrl_inst.latch_mem_inst.gclk\[8\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[8\]\[7\] sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_24_311 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_447 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_347 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[19\].gen_latches\[6\].p_latch net193 dig_ctrl_inst.latch_mem_inst.gclk\[19\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[19\]\[6\] sky130_fd_sc_hd__dlxtp_1
X_2483_ clknet_leaf_3_clk net336 net173 VGND VGND VDPWR VDPWR dig_ctrl_inst.spi_receiver_inst.spi_mosi_sync
+ sky130_fd_sc_hd__dfrtp_1
X_1503_ _1004_ _0211_ _0218_ _0204_ VGND VGND VDPWR VDPWR _0022_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_2_324 VDPWR VGND VDPWR VGND sky130_ef_sc_hd__decap_12
X_1434_ net251 _1039_ net15 VGND VGND VDPWR VDPWR net27 sky130_fd_sc_hd__mux2_1
X_1365_ net107 net101 net59 VGND VGND VDPWR VDPWR _0139_ sky130_fd_sc_hd__and3_2
X_1296_ _1075_ _1077_ _1093_ net135 net136 VGND VGND VDPWR VDPWR _1138_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_5_195 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_135 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_44_428 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_27 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_1150_ dig_ctrl_inst.cpu_inst.cpu_state\[2\] VGND VGND VDPWR VDPWR _0999_ sky130_fd_sc_hd__inv_2
XFILLER_0_23_42 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_8
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[5\].clock_gate clknet_leaf_0_clk dig_ctrl_inst.latch_mem_inst.data_we\[5\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.gen_gclk\[5\]._gclk sky130_fd_sc_hd__dlclkp_1
XFILLER_0_55_341 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_1983_ dig_ctrl_inst.latch_mem_inst.RAM\[50\]\[7\] net110 net47 VGND VGND VDPWR VDPWR
+ _0688_ sky130_fd_sc_hd__and3_2
X_1417_ net250 dig_ctrl_inst.spi_data_o\[2\] _1054_ _0162_ VGND VGND VDPWR VDPWR dig_ctrl_inst.data_out\[2\]
+ sky130_fd_sc_hd__a22o_1
X_2466_ clknet_leaf_7_clk _0072_ net143 VGND VGND VDPWR VDPWR dig_ctrl_inst.cpu_inst.r3\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_1348_ net153 _0131_ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.data_we\[29\]
+ sky130_fd_sc_hd__and2_1
X_2397_ clknet_leaf_2_clk _0006_ net172 VGND VGND VDPWR VDPWR dig_ctrl_inst.spi_addr\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_1279_ _1113_ _1120_ _1126_ dig_ctrl_inst.spi_addr\[4\] _1002_ VGND VGND VDPWR VDPWR
+ _1127_ sky130_fd_sc_hd__o32a_4
XTAP_TAPCELL_ROW_41_409 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout173 net176 VGND VGND VDPWR VDPWR net173 sky130_fd_sc_hd__clkbuf_4
Xfanout195 net196 VGND VGND VDPWR VDPWR net195 sky130_fd_sc_hd__clkbuf_2
Xfanout162 _1090_ VGND VGND VDPWR VDPWR net162 sky130_fd_sc_hd__buf_1
Xfanout140 net147 VGND VGND VDPWR VDPWR net140 sky130_fd_sc_hd__clkbuf_4
Xfanout151 net152 VGND VGND VDPWR VDPWR net151 sky130_fd_sc_hd__clkbuf_2
Xfanout184 net190 VGND VGND VDPWR VDPWR net184 sky130_fd_sc_hd__buf_2
XFILLER_0_56_149 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_341 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_2320_ dig_ctrl_inst.spi_receiver_inst.spi_cnt\[1\] _0980_ VGND VGND VDPWR VDPWR
+ _0981_ sky130_fd_sc_hd__and2b_1
XFILLER_0_69_49 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_2251_ _0229_ _0785_ _0792_ _0228_ VGND VGND VDPWR VDPWR _0938_ sky130_fd_sc_hd__a2bb2o_1
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[53\].clock_buffer dig_ctrl_inst.latch_mem_inst.gen_gclk\[53\]._gclk
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.gclk\[53\] sky130_fd_sc_hd__clkbuf_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[52\].gen_latches\[6\].p_latch net191 dig_ctrl_inst.latch_mem_inst.gclk\[52\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[52\]\[6\] sky130_fd_sc_hd__dlxtp_1
X_1202_ net260 net256 dig_ctrl_inst.cpu_inst.r2\[2\] VGND VGND VDPWR VDPWR _1050_
+ sky130_fd_sc_hd__and3b_1
X_2182_ _0252_ _0787_ _0825_ net166 VGND VGND VDPWR VDPWR _0872_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_18_97 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
X_1966_ dig_ctrl_inst.latch_mem_inst.RAM\[11\]\[6\] _1145_ _0637_ _0638_ _0649_ VGND
+ VGND VDPWR VDPWR _0672_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_63_545 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_40 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_41 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[41\].gen_latches\[4\].p_latch net210 dig_ctrl_inst.latch_mem_inst.gclk\[41\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[41\]\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_70_141 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[30\].gen_latches\[2\].p_latch net230 dig_ctrl_inst.latch_mem_inst.gclk\[30\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[30\]\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_55_182 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_95 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_1897_ dig_ctrl_inst.latch_mem_inst.RAM\[20\]\[5\] net98 net63 VGND VGND VDPWR VDPWR
+ _0604_ sky130_fd_sc_hd__and3_2
X_2449_ clknet_leaf_6_clk _0057_ net144 VGND VGND VDPWR VDPWR dig_ctrl_inst.cpu_inst.r1\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_2518_ clknet_leaf_11_clk VGND VGND VDPWR VDPWR net16 sky130_fd_sc_hd__buf_2
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[33\].clock_gate clknet_leaf_12_clk dig_ctrl_inst.latch_mem_inst.data_we\[33\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.gen_gclk\[33\]._gclk sky130_fd_sc_hd__dlclkp_1
XFILLER_0_19_341 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_77_626 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[56\].gen_latches\[7\].p_latch net188 dig_ctrl_inst.latch_mem_inst.gclk\[56\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[56\]\[7\] sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_60_526 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_160 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_17_269 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1820_ dig_ctrl_inst.latch_mem_inst.RAM\[48\]\[4\] net129 net45 VGND VGND VDPWR VDPWR
+ _0528_ sky130_fd_sc_hd__and3_2
X_1751_ dig_ctrl_inst.latch_mem_inst.RAM\[60\]\[3\] _0157_ _0278_ dig_ctrl_inst.latch_mem_inst.RAM\[5\]\[3\]
+ VGND VGND VDPWR VDPWR _0460_ sky130_fd_sc_hd__a22o_1
XFILLER_0_52_152 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_1682_ dig_ctrl_inst.latch_mem_inst.RAM\[17\]\[1\] _0120_ _0350_ _0358_ _0371_ VGND
+ VGND VDPWR VDPWR _0393_ sky130_fd_sc_hd__a2111o_1
Xmax_cap137 _0759_ VGND VGND VDPWR VDPWR net137 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_20_65 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_2303_ net381 _0971_ _0976_ VGND VGND VDPWR VDPWR _0064_ sky130_fd_sc_hd__mux2_1
X_2234_ _1110_ _0901_ VGND VGND VDPWR VDPWR _0922_ sky130_fd_sc_hd__xor2_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[45\].gen_latches\[5\].p_latch net199 dig_ctrl_inst.latch_mem_inst.gclk\[45\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[45\]\[5\] sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[1\].gen_latches\[0\].p_latch net240 dig_ctrl_inst.latch_mem_inst.gclk\[1\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[1\]\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_45_40 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_2165_ _1060_ _0829_ VGND VGND VDPWR VDPWR _0856_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_0_159 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2096_ _0787_ _0788_ _0261_ VGND VGND VDPWR VDPWR _0789_ sky130_fd_sc_hd__a21bo_1
X_1949_ dig_ctrl_inst.latch_mem_inst.RAM\[36\]\[6\] net97 net57 VGND VGND VDPWR VDPWR
+ _0655_ sky130_fd_sc_hd__and3_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[34\].gen_latches\[3\].p_latch net219 dig_ctrl_inst.latch_mem_inst.gclk\[34\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[34\]\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_0_53 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_75 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
X_2522__271 VGND VGND VDPWR VDPWR _2522__271/HI net271 sky130_fd_sc_hd__conb_1
XFILLER_0_43_196 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_8_215 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_74_607 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[23\].gen_latches\[1\].p_latch net238 dig_ctrl_inst.latch_mem_inst.gclk\[23\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[23\]\[1\] sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_22_294 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_13_Right_13 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_54 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_222 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
X_1803_ _0509_ _0510_ VGND VGND VDPWR VDPWR _0511_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_22_Right_22 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
X_1734_ dig_ctrl_inst.latch_mem_inst.RAM\[26\]\[2\] _0129_ _0156_ dig_ctrl_inst.latch_mem_inst.RAM\[59\]\[2\]
+ VGND VGND VDPWR VDPWR _0444_ sky130_fd_sc_hd__a22o_1
X_1596_ dig_ctrl_inst.latch_mem_inst.RAM\[3\]\[0\] _1135_ _0134_ dig_ctrl_inst.latch_mem_inst.RAM\[32\]\[0\]
+ _0307_ VGND VGND VDPWR VDPWR _0308_ sky130_fd_sc_hd__a221o_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[5\].gen_latches\[1\].p_latch net237 dig_ctrl_inst.latch_mem_inst.gclk\[5\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[5\]\[1\] sky130_fd_sc_hd__dlxtp_1
X_1665_ dig_ctrl_inst.latch_mem_inst.RAM\[54\]\[1\] _0152_ _0160_ dig_ctrl_inst.latch_mem_inst.RAM\[63\]\[1\]
+ _0375_ VGND VGND VDPWR VDPWR _0376_ sky130_fd_sc_hd__a221o_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[49\].gen_latches\[6\].p_latch net197 dig_ctrl_inst.latch_mem_inst.gclk\[49\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[49\]\[6\] sky130_fd_sc_hd__dlxtp_1
X_2217_ _0900_ _0905_ _0883_ VGND VGND VDPWR VDPWR _0049_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_31_Right_31 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_3 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[38\].gen_latches\[4\].p_latch net213 dig_ctrl_inst.latch_mem_inst.gclk\[38\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[38\]\[4\] sky130_fd_sc_hd__dlxtp_1
X_2148_ _0763_ _0768_ _0777_ _0765_ _0772_ VGND VGND VDPWR VDPWR _0839_ sky130_fd_sc_hd__o221a_1
X_2079_ net168 _0764_ VGND VGND VDPWR VDPWR _0772_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_40_Right_40 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_111 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_155 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[27\].gen_latches\[2\].p_latch net227 dig_ctrl_inst.latch_mem_inst.gclk\[27\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[27\]\[2\] sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[16\].gen_latches\[0\].p_latch net240 dig_ctrl_inst.latch_mem_inst.gclk\[16\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[16\]\[0\] sky130_fd_sc_hd__dlxtp_1
X_1450_ net391 _0182_ VGND VGND VDPWR VDPWR _0004_ sky130_fd_sc_hd__xor2_1
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[46\].clock_buffer dig_ctrl_inst.latch_mem_inst.gen_gclk\[46\]._gclk
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.gclk\[46\] sky130_fd_sc_hd__clkbuf_4
X_1381_ net152 _0146_ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.data_we\[47\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_77_306 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
X_2002_ dig_ctrl_inst.latch_mem_inst.RAM\[2\]\[7\] net121 net111 VGND VGND VDPWR VDPWR
+ _0707_ sky130_fd_sc_hd__and3_2
XFILLER_0_45_225 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[9\].gen_latches\[2\].p_latch net228 dig_ctrl_inst.latch_mem_inst.gclk\[9\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[9\]\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_5_322 VDPWR VGND VDPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_155 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
X_1648_ dig_ctrl_inst.latch_mem_inst.RAM\[40\]\[1\] net86 net52 VGND VGND VDPWR VDPWR
+ _0359_ sky130_fd_sc_hd__and3_2
X_1579_ dig_ctrl_inst.latch_mem_inst.RAM\[1\]\[0\] net131 net122 net116 VGND VGND
+ VDPWR VDPWR _0291_ sky130_fd_sc_hd__and4_1
X_1717_ dig_ctrl_inst.latch_mem_inst.RAM\[3\]\[2\] _1135_ _0157_ dig_ctrl_inst.latch_mem_inst.RAM\[60\]\[2\]
+ _0424_ VGND VGND VDPWR VDPWR _0427_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_16_Left_94 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_182 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_55_492 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_448 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_228 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
X_2482_ clknet_leaf_3_clk net12 net173 VGND VGND VDPWR VDPWR dig_ctrl_inst.spi_receiver_inst.synchronizer_spi_mosi.pipe\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_1433_ dig_ctrl_inst.port_ms_sync_i dig_ctrl_inst.spi_receiver_inst.stb_o net15 VGND
+ VGND VDPWR VDPWR net26 sky130_fd_sc_hd__mux2_1
X_1502_ _0174_ _0217_ _0216_ VGND VGND VDPWR VDPWR _0218_ sky130_fd_sc_hd__o21a_1
XFILLER_0_2_336 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_103 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
X_1295_ net153 net124 net118 _1136_ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.data_we\[5\]
+ sky130_fd_sc_hd__and4_1
X_1364_ net149 net93 net51 VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.data_we\[38\]
+ sky130_fd_sc_hd__and3_2
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[38\].clock_gate clknet_leaf_17_clk dig_ctrl_inst.latch_mem_inst.data_we\[38\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.gen_gclk\[38\]._gclk sky130_fd_sc_hd__dlclkp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[60\].gen_latches\[2\].p_latch net224 dig_ctrl_inst.latch_mem_inst.gclk\[60\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[60\]\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_68_125 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_44_429 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_1_Left_79 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[3\].clock_buffer dig_ctrl_inst.latch_mem_inst.gen_gclk\[3\]._gclk
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.gclk\[3\] sky130_fd_sc_hd__clkbuf_4
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[40\].clock_gate clknet_leaf_17_clk dig_ctrl_inst.latch_mem_inst.data_we\[40\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.gen_gclk\[40\]._gclk sky130_fd_sc_hd__dlclkp_1
XFILLER_0_59_169 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
X_1982_ dig_ctrl_inst.latch_mem_inst.RAM\[45\]\[7\] net115 net80 net52 VGND VGND VDPWR
+ VDPWR _0687_ sky130_fd_sc_hd__and4_1
XFILLER_0_30_209 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
X_1347_ net118 net82 net70 VGND VGND VDPWR VDPWR _0131_ sky130_fd_sc_hd__and3_2
X_2396_ clknet_leaf_3_clk _0005_ net172 VGND VGND VDPWR VDPWR dig_ctrl_inst.spi_addr\[0\]
+ sky130_fd_sc_hd__dfrtp_2
X_1416_ net250 dig_ctrl_inst.spi_data_o\[1\] _1084_ _0162_ VGND VGND VDPWR VDPWR dig_ctrl_inst.data_out\[1\]
+ sky130_fd_sc_hd__a22o_1
X_2465_ clknet_leaf_8_clk _0071_ net143 VGND VGND VDPWR VDPWR dig_ctrl_inst.cpu_inst.r3\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_64_94 VDPWR VGND VDPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_83 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_1278_ _1039_ _1125_ net249 VGND VGND VDPWR VDPWR _1126_ sky130_fd_sc_hd__a21o_1
XFILLER_0_3_42 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
XFILLER_0_65_139 VDPWR VGND VDPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_106 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_6
X_2525__280 VGND VGND VDPWR VDPWR net280 _2525__280/LO sky130_fd_sc_hd__conb_1
XFILLER_0_14_250 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
Xfanout174 net176 VGND VGND VDPWR VDPWR net174 sky130_fd_sc_hd__clkbuf_4
Xfanout196 net198 VGND VGND VDPWR VDPWR net196 sky130_fd_sc_hd__buf_1
Xfanout130 _1095_ VGND VGND VDPWR VDPWR net130 sky130_fd_sc_hd__buf_2
Xfanout185 net186 VGND VGND VDPWR VDPWR net185 sky130_fd_sc_hd__clkbuf_2
Xfanout141 net142 VGND VGND VDPWR VDPWR net141 sky130_fd_sc_hd__clkbuf_4
Xfanout152 _1097_ VGND VGND VDPWR VDPWR net152 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_6_198 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout163 _1084_ VGND VGND VDPWR VDPWR net163 sky130_fd_sc_hd__buf_8
XPHY_EDGE_ROW_69_Right_69 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[53\].gen_latches\[1\].p_latch net234 dig_ctrl_inst.latch_mem_inst.gclk\[53\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[53\]\[1\] sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[39\].clock_buffer dig_ctrl_inst.latch_mem_inst.gen_gclk\[39\]._gclk
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.gclk\[39\] sky130_fd_sc_hd__clkbuf_4
X_1201_ net182 net297 _1027_ dig_ctrl_inst.cpu_inst.ip\[2\] VGND VGND VDPWR VDPWR
+ _1049_ sky130_fd_sc_hd__o211a_1
X_2250_ dig_ctrl_inst.cpu_inst.data\[6\] _0743_ _0825_ net160 VGND VGND VDPWR VDPWR
+ _0937_ sky130_fd_sc_hd__a22o_1
XFILLER_0_34_64 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
X_2181_ net170 _0786_ _0793_ _0249_ VGND VGND VDPWR VDPWR _0871_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_71_590 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1965_ _0667_ _0668_ _0669_ _0670_ VGND VGND VDPWR VDPWR _0671_ sky130_fd_sc_hd__or4_1
X_2517_ clknet_leaf_3_clk net251 net173 VGND VGND VDPWR VDPWR dig_ctrl_inst.mode_d
+ sky130_fd_sc_hd__dfrtp_1
X_1896_ _0599_ _0600_ _0601_ _0602_ VGND VGND VDPWR VDPWR _0603_ sky130_fd_sc_hd__or4_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[30\].gen_latches\[6\].p_latch net195 dig_ctrl_inst.latch_mem_inst.gclk\[30\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[30\]\[6\] sky130_fd_sc_hd__dlxtp_1
X_2379_ clknet_leaf_4_clk net339 net174 VGND VGND VDPWR VDPWR dig_ctrl_inst.synchronizer_port_i_inst\[7\].out
+ sky130_fd_sc_hd__dfrtp_1
X_2448_ clknet_leaf_6_clk _0056_ net145 VGND VGND VDPWR VDPWR dig_ctrl_inst.cpu_inst.r1\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_52_3 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_139 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_194 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_183 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_77_627 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[57\].gen_latches\[2\].p_latch net224 dig_ctrl_inst.latch_mem_inst.gclk\[57\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[57\]\[2\] sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_60_527 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1750_ _0287_ _0451_ _0453_ _0458_ VGND VGND VDPWR VDPWR _0459_ sky130_fd_sc_hd__nor4_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[46\].gen_latches\[0\].p_latch net245 dig_ctrl_inst.latch_mem_inst.gclk\[46\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[46\]\[0\] sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_4_Left_82 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_315 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_6
X_1681_ dig_ctrl_inst.latch_mem_inst.RAM\[45\]\[1\] _0145_ _0348_ _0365_ _0370_ VGND
+ VGND VDPWR VDPWR _0392_ sky130_fd_sc_hd__a2111o_1
X_2164_ dig_ctrl_inst.synchronizer_port_i_inst\[2\].out _0802_ _0804_ dig_ctrl_inst.spi_data_o\[2\]
+ VGND VGND VDPWR VDPWR _0855_ sky130_fd_sc_hd__a22oi_1
X_2302_ net371 _0970_ _0976_ VGND VGND VDPWR VDPWR _0063_ sky130_fd_sc_hd__mux2_1
X_2233_ _1110_ _1125_ _0878_ VGND VGND VDPWR VDPWR _0921_ sky130_fd_sc_hd__and3_2
XFILLER_0_29_53 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[1\].gen_latches\[4\].p_latch net214 dig_ctrl_inst.latch_mem_inst.gclk\[1\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[1\]\[4\] sky130_fd_sc_hd__dlxtp_1
X_2095_ _1014_ _0744_ VGND VGND VDPWR VDPWR _0788_ sky130_fd_sc_hd__or2_4
X_1948_ dig_ctrl_inst.latch_mem_inst.RAM\[47\]\[6\] net107 _1146_ net57 VGND VGND
+ VDPWR VDPWR _0654_ sky130_fd_sc_hd__and4_1
XFILLER_0_9_63 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_1879_ dig_ctrl_inst.latch_mem_inst.RAM\[35\]\[5\] _0137_ _0583_ _0584_ _0585_ VGND
+ VGND VDPWR VDPWR _0586_ sky130_fd_sc_hd__a2111o_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[34\].gen_latches\[7\].p_latch net185 dig_ctrl_inst.latch_mem_inst.gclk\[34\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[34\]\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_31_337 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_74_608 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[10\].clock_buffer dig_ctrl_inst.latch_mem_inst.gen_gclk\[10\]._gclk
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.gclk\[10\] sky130_fd_sc_hd__clkbuf_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[23\].gen_latches\[5\].p_latch net201 dig_ctrl_inst.latch_mem_inst.gclk\[23\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[23\]\[5\] sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[12\].gen_latches\[3\].p_latch net222 dig_ctrl_inst.latch_mem_inst.gclk\[12\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[12\]\[3\] sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_22_295 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_29 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_1802_ dig_ctrl_inst.latch_mem_inst.RAM\[50\]\[4\] net110 net44 _1133_ dig_ctrl_inst.latch_mem_inst.RAM\[2\]\[4\]
+ VGND VGND VDPWR VDPWR _0510_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_13_240 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1733_ dig_ctrl_inst.latch_mem_inst.RAM\[25\]\[2\] _0128_ _0154_ dig_ctrl_inst.latch_mem_inst.RAM\[57\]\[2\]
+ VGND VGND VDPWR VDPWR _0443_ sky130_fd_sc_hd__a22o_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[5\].gen_latches\[5\].p_latch net205 dig_ctrl_inst.latch_mem_inst.gclk\[5\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[5\]\[5\] sky130_fd_sc_hd__dlxtp_1
X_1595_ dig_ctrl_inst.latch_mem_inst.RAM\[40\]\[0\] _0140_ _0156_ dig_ctrl_inst.latch_mem_inst.RAM\[59\]\[0\]
+ VGND VGND VDPWR VDPWR _0307_ sky130_fd_sc_hd__a22o_1
X_1664_ dig_ctrl_inst.latch_mem_inst.RAM\[56\]\[1\] net88 net50 _0131_ dig_ctrl_inst.latch_mem_inst.RAM\[29\]\[1\]
+ VGND VGND VDPWR VDPWR _0375_ sky130_fd_sc_hd__a32o_1
XFILLER_0_0_253 VDPWR VGND VDPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_337 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
X_2216_ _0754_ _0903_ _0904_ _0756_ net41 VGND VGND VDPWR VDPWR _0905_ sky130_fd_sc_hd__o221a_1
X_2147_ _0264_ _0760_ _0836_ _0837_ _0770_ VGND VGND VDPWR VDPWR _0838_ sky130_fd_sc_hd__o32a_1
X_2078_ _0264_ _0760_ _0770_ VGND VGND VDPWR VDPWR _0771_ sky130_fd_sc_hd__or3_1
XFILLER_0_71_281 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_134 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_8
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[45\].clock_gate clknet_leaf_16_clk dig_ctrl_inst.latch_mem_inst.data_we\[45\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.gen_gclk\[45\]._gclk sky130_fd_sc_hd__dlclkp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[27\].gen_latches\[6\].p_latch net198 dig_ctrl_inst.latch_mem_inst.gclk\[27\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[27\]\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_39_223 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[16\].gen_latches\[4\].p_latch net208 dig_ctrl_inst.latch_mem_inst.gclk\[16\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[16\]\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_10_307 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_1380_ net104 net81 net54 VGND VGND VDPWR VDPWR _0146_ sky130_fd_sc_hd__and3_4
X_2001_ dig_ctrl_inst.latch_mem_inst.RAM\[61\]\[7\] net115 net80 net42 VGND VGND VDPWR
+ VDPWR _0706_ sky130_fd_sc_hd__and4_1
XFILLER_0_42_75 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_8
Xdig_ctrl_inst.latch_mem_inst.gen_words\[9\].gen_latches\[6\].p_latch net197 dig_ctrl_inst.latch_mem_inst.gclk\[9\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[9\]\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_5_334 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_167 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_1716_ dig_ctrl_inst.latch_mem_inst.RAM\[35\]\[2\] _0137_ _0145_ dig_ctrl_inst.latch_mem_inst.RAM\[45\]\[2\]
+ _0425_ VGND VGND VDPWR VDPWR _0426_ sky130_fd_sc_hd__a221o_1
X_1578_ dig_ctrl_inst.latch_mem_inst.RAM\[23\]\[0\] net108 net101 net71 VGND VGND
+ VDPWR VDPWR _0290_ sky130_fd_sc_hd__and4_1
X_1647_ dig_ctrl_inst.latch_mem_inst.RAM\[19\]\[1\] net133 net105 net66 VGND VGND
+ VDPWR VDPWR _0358_ sky130_fd_sc_hd__and4_1
Xrebuffer20 net303 VGND VGND VDPWR VDPWR net302 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_4_3 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_55_493 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_449 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2481_ clknet_leaf_3_clk net344 VGND VGND VDPWR VDPWR dig_ctrl_inst.spi_receiver_inst.spi_sclk_delayed
+ sky130_fd_sc_hd__dfxtp_1
X_1363_ net156 _0138_ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.data_we\[37\]
+ sky130_fd_sc_hd__and2_1
X_1432_ net250 dig_ctrl_inst.spi_data_o\[7\] _0162_ _0172_ VGND VGND VDPWR VDPWR dig_ctrl_inst.data_out\[7\]
+ sky130_fd_sc_hd__a22o_1
X_1501_ net169 dig_ctrl_inst.cpu_inst.data\[3\] _0198_ VGND VGND VDPWR VDPWR _0217_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_148 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
X_1294_ net154 net125 net97 VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.data_we\[4\]
+ sky130_fd_sc_hd__and3_2
XFILLER_0_53_41 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XFILLER_0_58_340 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[60\].gen_latches\[6\].p_latch net322 dig_ctrl_inst.latch_mem_inst.gclk\[60\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[60\]\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_64_321 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_52_474 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_281 VDPWR VGND VDPWR VGND sky130_ef_sc_hd__decap_12
X_1981_ dig_ctrl_inst.latch_mem_inst.RAM\[0\]\[7\] _0288_ VGND VGND VDPWR VDPWR _0686_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_15_229 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_6
X_1346_ net153 net78 net70 VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.data_we\[28\]
+ sky130_fd_sc_hd__and3_2
X_2395_ clknet_leaf_6_clk net340 net180 VGND VGND VDPWR VDPWR dig_ctrl_inst.port_ms_sync_i
+ sky130_fd_sc_hd__dfrtp_1
X_1415_ net250 dig_ctrl_inst.spi_data_o\[0\] _1067_ _0162_ VGND VGND VDPWR VDPWR dig_ctrl_inst.data_out\[0\]
+ sky130_fd_sc_hd__a22o_1
X_2464_ clknet_leaf_10_clk _0070_ net139 VGND VGND VDPWR VDPWR dig_ctrl_inst.cpu_inst.r3\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_64_51 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_1277_ _1021_ _1121_ _1122_ _1123_ _1124_ VGND VGND VDPWR VDPWR _1125_ sky130_fd_sc_hd__o41a_2
Xfanout120 net122 VGND VGND VDPWR VDPWR net120 sky130_fd_sc_hd__buf_2
Xfanout131 net133 VGND VGND VDPWR VDPWR net131 sky130_fd_sc_hd__buf_2
XFILLER_0_14_273 VDPWR VGND VDPWR VGND sky130_ef_sc_hd__decap_12
Xfanout175 net176 VGND VGND VDPWR VDPWR net175 sky130_fd_sc_hd__clkbuf_2
Xfanout153 net154 VGND VGND VDPWR VDPWR net153 sky130_fd_sc_hd__clkbuf_2
Xfanout197 net198 VGND VGND VDPWR VDPWR net197 sky130_fd_sc_hd__clkbuf_2
Xfanout186 net190 VGND VGND VDPWR VDPWR net186 sky130_fd_sc_hd__clkbuf_2
Xfanout142 net147 VGND VGND VDPWR VDPWR net142 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_6_199 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout164 net295 VGND VGND VDPWR VDPWR net164 sky130_fd_sc_hd__buf_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[53\].gen_latches\[5\].p_latch net199 dig_ctrl_inst.latch_mem_inst.gclk\[53\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[53\]\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_69_18 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[42\].gen_latches\[3\].p_latch net222 dig_ctrl_inst.latch_mem_inst.gclk\[42\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[42\]\[3\] sky130_fd_sc_hd__dlxtp_1
X_1200_ net249 _1029_ _1046_ _1038_ _1008_ VGND VGND VDPWR VDPWR _1048_ sky130_fd_sc_hd__o41ai_4
XFILLER_0_18_33 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_2180_ dig_ctrl_inst.cpu_inst.data\[3\] _0743_ _0785_ _0250_ VGND VGND VDPWR VDPWR
+ _0870_ sky130_fd_sc_hd__o2bb2a_1
XTAP_TAPCELL_ROW_71_591 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1964_ dig_ctrl_inst.latch_mem_inst.RAM\[29\]\[6\] _0131_ _0144_ dig_ctrl_inst.latch_mem_inst.RAM\[44\]\[6\]
+ _0662_ VGND VGND VDPWR VDPWR _0670_ sky130_fd_sc_hd__a221o_1
X_1895_ dig_ctrl_inst.latch_mem_inst.RAM\[47\]\[5\] _0146_ _0160_ dig_ctrl_inst.latch_mem_inst.RAM\[63\]\[5\]
+ VGND VGND VDPWR VDPWR _0602_ sky130_fd_sc_hd__a22o_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[31\].gen_latches\[1\].p_latch net233 dig_ctrl_inst.latch_mem_inst.gclk\[31\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[31\]\[1\] sky130_fd_sc_hd__dlxtp_1
Xclkbuf_leaf_13_clk clknet_1_0__leaf_clk VGND VGND VDPWR VDPWR clknet_leaf_13_clk
+ sky130_fd_sc_hd__clkbuf_8
X_2447_ clknet_leaf_8_clk _0055_ net146 VGND VGND VDPWR VDPWR dig_ctrl_inst.cpu_inst.r1\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_2516_ clknet_leaf_8_clk _0113_ net143 VGND VGND VDPWR VDPWR dig_ctrl_inst.cpu_inst.cpu_state\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_2378_ clknet_leaf_3_clk net10 net173 VGND VGND VDPWR VDPWR dig_ctrl_inst.synchronizer_port_i_inst\[7\].pipe\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_1329_ net154 _0122_ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.data_we\[19\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_45_3 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_77_628 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[57\].gen_latches\[6\].p_latch net194 dig_ctrl_inst.latch_mem_inst.gclk\[57\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[57\]\[6\] sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[52\].clock_gate clknet_leaf_12_clk dig_ctrl_inst.latch_mem_inst.data_we\[52\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.gen_gclk\[52\]._gclk sky130_fd_sc_hd__dlclkp_1
X_2301_ net362 _0969_ _0976_ VGND VGND VDPWR VDPWR _0062_ sky130_fd_sc_hd__mux2_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[46\].gen_latches\[4\].p_latch net210 dig_ctrl_inst.latch_mem_inst.gclk\[46\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[46\]\[4\] sky130_fd_sc_hd__dlxtp_1
X_1680_ _0387_ _0388_ _0389_ _0390_ VGND VGND VDPWR VDPWR _0391_ sky130_fd_sc_hd__or4_1
Xclkbuf_leaf_2_clk clknet_1_1__leaf_clk VGND VGND VDPWR VDPWR clknet_leaf_2_clk sky130_fd_sc_hd__clkbuf_8
X_2163_ _0788_ _0853_ _0851_ _0841_ VGND VGND VDPWR VDPWR _0854_ sky130_fd_sc_hd__o211a_1
X_2232_ _0788_ _0907_ _0910_ _0919_ VGND VGND VDPWR VDPWR _0920_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_61_63 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_2094_ _0742_ _0745_ VGND VGND VDPWR VDPWR _0787_ sky130_fd_sc_hd__or2_2
XTAP_TAPCELL_ROW_16_260 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[35\].gen_latches\[2\].p_latch net224 dig_ctrl_inst.latch_mem_inst.gclk\[35\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[35\]\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_43_143 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_195 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_1878_ dig_ctrl_inst.latch_mem_inst.RAM\[31\]\[5\] net102 net81 net62 VGND VGND VDPWR
+ VDPWR _0585_ sky130_fd_sc_hd__and4_1
XFILLER_0_9_53 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
X_1947_ dig_ctrl_inst.latch_mem_inst.RAM\[14\]\[6\] net120 net75 VGND VGND VDPWR VDPWR
+ _0653_ sky130_fd_sc_hd__and3_2
XFILLER_0_16_302 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[24\].gen_latches\[0\].p_latch net240 dig_ctrl_inst.latch_mem_inst.gclk\[24\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[24\]\[0\] sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_74_609 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_396 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_224 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_140 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_22_296 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[12\].gen_latches\[7\].p_latch net183 dig_ctrl_inst.latch_mem_inst.gclk\[12\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[12\]\[7\] sky130_fd_sc_hd__dlxtp_1
X_1732_ _0440_ _0441_ VGND VGND VDPWR VDPWR _0442_ sky130_fd_sc_hd__or2_1
X_1663_ dig_ctrl_inst.latch_mem_inst.RAM\[4\]\[1\] _0277_ _0278_ dig_ctrl_inst.latch_mem_inst.RAM\[5\]\[1\]
+ _0373_ VGND VGND VDPWR VDPWR _0374_ sky130_fd_sc_hd__a221o_1
XFILLER_0_40_124 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[6\].gen_latches\[0\].p_latch net241 dig_ctrl_inst.latch_mem_inst.gclk\[6\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[6\]\[0\] sky130_fd_sc_hd__dlxtp_1
X_1801_ dig_ctrl_inst.latch_mem_inst.RAM\[46\]\[4\] net75 net55 _0137_ dig_ctrl_inst.latch_mem_inst.RAM\[35\]\[4\]
+ VGND VGND VDPWR VDPWR _0509_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_13_241 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_316 VDPWR VGND VDPWR VGND sky130_ef_sc_hd__decap_12
X_1594_ dig_ctrl_inst.latch_mem_inst.RAM\[2\]\[0\] _1133_ _0139_ dig_ctrl_inst.latch_mem_inst.RAM\[39\]\[0\]
+ _0305_ VGND VGND VDPWR VDPWR _0306_ sky130_fd_sc_hd__a221o_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[39\].gen_latches\[3\].p_latch net218 dig_ctrl_inst.latch_mem_inst.gclk\[39\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[39\]\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_0_265 VDPWR VGND VDPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_7_Right_7 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
X_2215_ dig_ctrl_inst.synchronizer_port_i_inst\[4\].out _0802_ _0804_ dig_ctrl_inst.spi_data_o\[4\]
+ VGND VGND VDPWR VDPWR _0904_ sky130_fd_sc_hd__a22oi_1
X_2146_ _0762_ _0766_ net157 VGND VGND VDPWR VDPWR _0837_ sky130_fd_sc_hd__mux2_1
X_2077_ net163 _0769_ VGND VGND VDPWR VDPWR _0770_ sky130_fd_sc_hd__nand2b_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[28\].gen_latches\[1\].p_latch net236 dig_ctrl_inst.latch_mem_inst.gclk\[28\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[28\]\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_31_113 VDPWR VGND VDPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_24_Left_102 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_33_Left_111 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_10_222 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_42_Left_120 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
X_2000_ dig_ctrl_inst.latch_mem_inst.RAM\[41\]\[7\] net114 net90 net51 VGND VGND VDPWR
+ VDPWR _0705_ sky130_fd_sc_hd__and4_1
X_1646_ dig_ctrl_inst.latch_mem_inst.RAM\[25\]\[1\] net115 net90 net61 VGND VGND VDPWR
+ VDPWR _0357_ sky130_fd_sc_hd__and4_1
X_1715_ dig_ctrl_inst.latch_mem_inst.RAM\[32\]\[2\] _0134_ _0158_ dig_ctrl_inst.latch_mem_inst.RAM\[61\]\[2\]
+ VGND VGND VDPWR VDPWR _0425_ sky130_fd_sc_hd__a22o_1
X_1577_ dig_ctrl_inst.latch_mem_inst.RAM\[34\]\[0\] net111 net58 VGND VGND VDPWR VDPWR
+ _0289_ sky130_fd_sc_hd__and3_2
XFILLER_0_6_98 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
Xrebuffer21 _1076_ VGND VGND VDPWR VDPWR net303 sky130_fd_sc_hd__clkbuf_1
Xrebuffer10 _1026_ VGND VGND VDPWR VDPWR net292 sky130_fd_sc_hd__dlygate4sd1_1
X_2129_ _0257_ _0258_ _0788_ VGND VGND VDPWR VDPWR _0821_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_36_249 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_195 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_55_494 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2480_ clknet_leaf_2_clk _0086_ net180 VGND VGND VDPWR VDPWR dig_ctrl_inst.spi_data_o\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_50_230 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
X_1500_ _0174_ _0215_ VGND VGND VDPWR VDPWR _0216_ sky130_fd_sc_hd__nand2_1
X_1293_ _1075_ _1077_ net134 net135 net136 VGND VGND VDPWR VDPWR _1137_ sky130_fd_sc_hd__o2111a_1
X_1362_ net118 net101 net57 VGND VGND VDPWR VDPWR _0138_ sky130_fd_sc_hd__and3_2
X_1431_ _1018_ _0168_ _0169_ _0170_ _0171_ VGND VGND VDPWR VDPWR _0172_ sky130_fd_sc_hd__o41a_4
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[42\].clock_buffer dig_ctrl_inst.latch_mem_inst.gen_gclk\[42\]._gclk
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.gclk\[42\] sky130_fd_sc_hd__clkbuf_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[61\].gen_latches\[1\].p_latch net232 dig_ctrl_inst.latch_mem_inst.gclk\[61\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[61\]\[1\] sky130_fd_sc_hd__dlxtp_1
X_1629_ dig_ctrl_inst.latch_mem_inst.RAM\[60\]\[1\] net76 net47 VGND VGND VDPWR VDPWR
+ _0340_ sky130_fd_sc_hd__and3_2
XTAP_TAPCELL_ROW_52_475 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[57\].clock_gate clknet_leaf_16_clk dig_ctrl_inst.latch_mem_inst.data_we\[57\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.gen_gclk\[57\]._gclk sky130_fd_sc_hd__dlclkp_1
XFILLER_0_17_271 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_293 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_105 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_43_420 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1980_ dig_ctrl_inst.cpu_inst.instr\[6\] _0685_ _0276_ VGND VGND VDPWR VDPWR _0032_
+ sky130_fd_sc_hd__mux2_1
X_2532_ net278 VGND VGND VDPWR VDPWR uio_out[5] sky130_fd_sc_hd__buf_2
Xrebuffer1 _1017_ VGND VGND VDPWR VDPWR net283 sky130_fd_sc_hd__buf_6
X_2463_ clknet_leaf_11_clk _0069_ net140 VGND VGND VDPWR VDPWR dig_ctrl_inst.cpu_inst.r3\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_1345_ net155 _0130_ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.data_we\[27\]
+ sky130_fd_sc_hd__and2_1
X_2394_ clknet_leaf_6_clk net1 net180 VGND VGND VDPWR VDPWR dig_ctrl_inst.synchronizer_port_ms_i_inst.pipe\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_1414_ net250 _1040_ VGND VGND VDPWR VDPWR _0162_ sky130_fd_sc_hd__nor2_2
XFILLER_0_48_97 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
X_1276_ net268 net263 dig_ctrl_inst.cpu_inst.r0\[4\] VGND VGND VDPWR VDPWR _1124_
+ sky130_fd_sc_hd__or3_1
XFILLER_0_3_11 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
Xfanout154 net155 VGND VGND VDPWR VDPWR net154 sky130_fd_sc_hd__clkbuf_2
Xfanout132 net133 VGND VGND VDPWR VDPWR net132 sky130_fd_sc_hd__clkbuf_4
Xfanout143 net147 VGND VGND VDPWR VDPWR net143 sky130_fd_sc_hd__clkbuf_4
Xfanout121 net122 VGND VGND VDPWR VDPWR net121 sky130_fd_sc_hd__clkbuf_2
Xfanout165 _1073_ VGND VGND VDPWR VDPWR net165 sky130_fd_sc_hd__buf_6
Xfanout110 net112 VGND VGND VDPWR VDPWR net110 sky130_fd_sc_hd__buf_2
XFILLER_0_14_285 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_6
Xdig_ctrl_inst.latch_mem_inst.gen_words\[54\].gen_latches\[0\].p_latch net240 dig_ctrl_inst.latch_mem_inst.gclk\[54\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[54\]\[0\] sky130_fd_sc_hd__dlxtp_1
Xfanout176 dig_ctrl_inst.latch_mem_inst.rst_ni VGND VGND VDPWR VDPWR net176 sky130_fd_sc_hd__clkbuf_2
Xfanout187 net188 VGND VGND VDPWR VDPWR net187 sky130_fd_sc_hd__buf_2
Xfanout198 net322 VGND VGND VDPWR VDPWR net198 sky130_fd_sc_hd__buf_2
XFILLER_0_64_141 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_160 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[42\].gen_latches\[7\].p_latch net188 dig_ctrl_inst.latch_mem_inst.gclk\[42\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[42\]\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_18_23 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_71_592 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_21 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_1963_ dig_ctrl_inst.latch_mem_inst.RAM\[20\]\[6\] _0123_ _0278_ dig_ctrl_inst.latch_mem_inst.RAM\[5\]\[6\]
+ _0661_ VGND VGND VDPWR VDPWR _0669_ sky130_fd_sc_hd__a221o_1
X_1894_ dig_ctrl_inst.latch_mem_inst.RAM\[50\]\[5\] net111 net45 _0138_ dig_ctrl_inst.latch_mem_inst.RAM\[37\]\[5\]
+ VGND VGND VDPWR VDPWR _0601_ sky130_fd_sc_hd__a32o_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[31\].gen_latches\[5\].p_latch net199 dig_ctrl_inst.latch_mem_inst.gclk\[31\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[31\]\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_59_41 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_2515_ clknet_leaf_9_clk _0112_ net142 VGND VGND VDPWR VDPWR dig_ctrl_inst.cpu_inst.cpu_state\[1\]
+ sky130_fd_sc_hd__dfrtp_4
X_2446_ clknet_leaf_9_clk _0054_ net141 VGND VGND VDPWR VDPWR dig_ctrl_inst.cpu_inst.r1\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_11_255 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_2377_ clknet_leaf_4_clk _0004_ net177 VGND VGND VDPWR VDPWR dig_ctrl_inst.spi_receiver_inst.spi_cnt\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_1328_ net132 net107 net70 VGND VGND VDPWR VDPWR _0122_ sky130_fd_sc_hd__and3_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[20\].gen_latches\[3\].p_latch net220 dig_ctrl_inst.latch_mem_inst.gclk\[20\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[20\]\[3\] sky130_fd_sc_hd__dlxtp_1
X_1259_ net267 net263 dig_ctrl_inst.cpu_inst.r3\[5\] VGND VGND VDPWR VDPWR _1107_
+ sky130_fd_sc_hd__and3_2
XFILLER_0_38_3 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_141 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_19_280 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_333 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_122 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[58\].gen_latches\[1\].p_latch net238 dig_ctrl_inst.latch_mem_inst.gclk\[58\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[58\]\[1\] sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_77_629 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_122 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[2\].gen_latches\[3\].p_latch net215 dig_ctrl_inst.latch_mem_inst.gclk\[2\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[2\]\[3\] sky130_fd_sc_hd__dlxtp_1
X_2231_ _0750_ _0912_ _0917_ _0918_ VGND VGND VDPWR VDPWR _0919_ sky130_fd_sc_hd__o211a_1
X_2300_ net379 _0968_ _0976_ VGND VGND VDPWR VDPWR _0061_ sky130_fd_sc_hd__mux2_1
XFILLER_0_45_54 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
X_2162_ _0248_ _0852_ VGND VGND VDPWR VDPWR _0853_ sky130_fd_sc_hd__xnor2_1
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[35\].clock_buffer dig_ctrl_inst.latch_mem_inst.gen_gclk\[35\]._gclk
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.gclk\[35\] sky130_fd_sc_hd__clkbuf_4
X_2093_ net253 _0745_ net252 VGND VGND VDPWR VDPWR _0786_ sky130_fd_sc_hd__or3b_4
XFILLER_0_75_225 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_163 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_16_261 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[35\].gen_latches\[6\].p_latch net194 dig_ctrl_inst.latch_mem_inst.gclk\[35\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[35\]\[6\] sky130_fd_sc_hd__dlxtp_1
X_1946_ dig_ctrl_inst.latch_mem_inst.RAM\[38\]\[6\] net95 net57 VGND VGND VDPWR VDPWR
+ _0652_ sky130_fd_sc_hd__and3_2
XFILLER_0_43_122 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
X_1877_ dig_ctrl_inst.latch_mem_inst.RAM\[53\]\[5\] net114 net99 net44 VGND VGND VDPWR
+ VDPWR _0584_ sky130_fd_sc_hd__and4_1
XFILLER_0_9_76 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[24\].gen_latches\[4\].p_latch net211 dig_ctrl_inst.latch_mem_inst.gclk\[24\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[24\]\[4\] sky130_fd_sc_hd__dlxtp_1
X_2429_ clknet_leaf_9_clk _0037_ net141 VGND VGND VDPWR VDPWR dig_ctrl_inst.cpu_inst.data\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_39_397 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[13\].gen_latches\[2\].p_latch net229 dig_ctrl_inst.latch_mem_inst.gclk\[13\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[13\]\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_34_166 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_111 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_22_297 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_203 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_1800_ dig_ctrl_inst.latch_mem_inst.RAM\[23\]\[4\] _0126_ _0279_ dig_ctrl_inst.latch_mem_inst.RAM\[6\]\[4\]
+ _0507_ VGND VGND VDPWR VDPWR _0508_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_13_242 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_57 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_1662_ dig_ctrl_inst.latch_mem_inst.RAM\[42\]\[1\] _0142_ _0148_ dig_ctrl_inst.latch_mem_inst.RAM\[49\]\[1\]
+ VGND VGND VDPWR VDPWR _0373_ sky130_fd_sc_hd__a22o_1
X_1731_ dig_ctrl_inst.latch_mem_inst.RAM\[46\]\[2\] net73 net57 _0138_ dig_ctrl_inst.latch_mem_inst.RAM\[37\]\[2\]
+ VGND VGND VDPWR VDPWR _0441_ sky130_fd_sc_hd__a32o_1
Xwire182 _1009_ VGND VGND VDPWR VDPWR net182 sky130_fd_sc_hd__clkbuf_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[6\].gen_latches\[4\].p_latch net211 dig_ctrl_inst.latch_mem_inst.gclk\[6\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[6\]\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_13_328 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_8
X_2214_ _0901_ _0902_ VGND VGND VDPWR VDPWR _0903_ sky130_fd_sc_hd__nand2_1
X_1593_ dig_ctrl_inst.latch_mem_inst.RAM\[20\]\[0\] _0123_ _0143_ dig_ctrl_inst.latch_mem_inst.RAM\[43\]\[0\]
+ VGND VGND VDPWR VDPWR _0305_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_277 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_97 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[39\].gen_latches\[7\].p_latch net189 dig_ctrl_inst.latch_mem_inst.gclk\[39\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[39\]\[7\] sky130_fd_sc_hd__dlxtp_1
X_2145_ net163 _0769_ VGND VGND VDPWR VDPWR _0836_ sky130_fd_sc_hd__nand2_2
X_2076_ net253 dig_ctrl_inst.cpu_inst.instr\[6\] dig_ctrl_inst.cpu_inst.instr\[7\]
+ net252 VGND VGND VDPWR VDPWR _0769_ sky130_fd_sc_hd__and4bb_1
XTAP_TAPCELL_ROW_36_378 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1929_ dig_ctrl_inst.latch_mem_inst.RAM\[24\]\[6\] net86 net64 VGND VGND VDPWR VDPWR
+ _0635_ sky130_fd_sc_hd__and3_2
XFILLER_0_16_166 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_169 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[28\].gen_latches\[5\].p_latch net202 dig_ctrl_inst.latch_mem_inst.gclk\[28\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[28\]\[5\] sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[17\].gen_latches\[3\].p_latch net217 dig_ctrl_inst.latch_mem_inst.gclk\[17\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[17\]\[3\] sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_10_223 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_309 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_6
Xhold90 net22 VGND VGND VDPWR VDPWR net372 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_5_314 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_272 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_1576_ _0284_ _0285_ _0286_ VGND VGND VDPWR VDPWR _0288_ sky130_fd_sc_hd__or3_4
XFILLER_0_6_11 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_1714_ dig_ctrl_inst.latch_mem_inst.RAM\[31\]\[2\] _0132_ _0135_ dig_ctrl_inst.latch_mem_inst.RAM\[33\]\[2\]
+ VGND VGND VDPWR VDPWR _0424_ sky130_fd_sc_hd__a22o_1
XFILLER_0_13_169 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
X_1645_ dig_ctrl_inst.latch_mem_inst.RAM\[14\]\[1\] net121 net72 VGND VGND VDPWR VDPWR
+ _0356_ sky130_fd_sc_hd__and3_2
XFILLER_0_67_52 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
Xrebuffer11 _1028_ VGND VGND VDPWR VDPWR net293 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_0_20_3 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
Xrebuffer22 _1076_ VGND VGND VDPWR VDPWR net304 sky130_fd_sc_hd__buf_2
X_2059_ _0751_ VGND VGND VDPWR VDPWR _0752_ sky130_fd_sc_hd__inv_2
X_2128_ net168 _0819_ _0813_ net171 VGND VGND VDPWR VDPWR _0820_ sky130_fd_sc_hd__a211o_1
XFILLER_0_12_180 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_55_495 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_209 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[28\].clock_buffer dig_ctrl_inst.latch_mem_inst.gen_gclk\[28\]._gclk
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.gclk\[28\] sky130_fd_sc_hd__clkbuf_4
X_1430_ net259 net254 dig_ctrl_inst.cpu_inst.r0\[7\] VGND VGND VDPWR VDPWR _0171_
+ sky130_fd_sc_hd__or3_1
XFILLER_0_10_139 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_1361_ net154 net97 net57 VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.data_we\[36\]
+ sky130_fd_sc_hd__and3_2
X_1292_ net136 net135 VGND VGND VDPWR VDPWR _1136_ sky130_fd_sc_hd__and2_4
XTAP_TAPCELL_ROW_46_440 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_3 VDPWR VGND VDPWR VGND sky130_ef_sc_hd__decap_12
Xdig_ctrl_inst.latch_mem_inst.gen_words\[61\].gen_latches\[5\].p_latch net199 dig_ctrl_inst.latch_mem_inst.gclk\[61\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[61\]\[5\] sky130_fd_sc_hd__dlxtp_1
X_1559_ _0237_ _0269_ _0270_ _0271_ net252 VGND VGND VDPWR VDPWR _0272_ sky130_fd_sc_hd__o2111ai_1
X_1628_ dig_ctrl_inst.latch_mem_inst.RAM\[39\]\[1\] net102 net99 net52 VGND VGND VDPWR
+ VDPWR _0339_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_69_576 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_61_Left_139 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XFILLER_0_68_139 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_52_476 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[50\].gen_latches\[3\].p_latch net215 dig_ctrl_inst.latch_mem_inst.gclk\[50\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[50\]\[3\] sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_70_Left_148 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_253 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_161 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_43_421 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer2 net283 VGND VGND VDPWR VDPWR net284 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_0_23_57 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
X_2462_ clknet_leaf_3_clk net335 net173 VGND VGND VDPWR VDPWR dig_ctrl_inst.mode_sync
+ sky130_fd_sc_hd__dfrtp_1
X_2531_ net277 VGND VGND VDPWR VDPWR uio_out[4] sky130_fd_sc_hd__buf_2
X_2393_ clknet_leaf_4_clk net341 net179 VGND VGND VDPWR VDPWR dig_ctrl_inst.synchronizer_port_i_inst\[0\].out
+ sky130_fd_sc_hd__dfrtp_1
X_1413_ _0161_ VGND VGND VDPWR VDPWR dig_ctrl_inst.cpu_inst.rst_ni sky130_fd_sc_hd__inv_2
XFILLER_0_2_147 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_125 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_253 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_1344_ net106 _1140_ net69 VGND VGND VDPWR VDPWR _0130_ sky130_fd_sc_hd__and3_2
XFILLER_0_64_20 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_1275_ net267 dig_ctrl_inst.cpu_inst.r2\[4\] VGND VGND VDPWR VDPWR _1123_ sky130_fd_sc_hd__and2b_1
XFILLER_0_3_23 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_337 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
Xfanout177 net180 VGND VGND VDPWR VDPWR net177 sky130_fd_sc_hd__clkbuf_4
Xfanout188 net189 VGND VGND VDPWR VDPWR net188 sky130_fd_sc_hd__buf_2
Xfanout133 _1063_ VGND VGND VDPWR VDPWR net133 sky130_fd_sc_hd__clkbuf_4
Xfanout155 net156 VGND VGND VDPWR VDPWR net155 sky130_fd_sc_hd__clkbuf_2
Xfanout111 net112 VGND VGND VDPWR VDPWR net111 sky130_fd_sc_hd__buf_2
Xfanout144 net147 VGND VGND VDPWR VDPWR net144 sky130_fd_sc_hd__clkbuf_2
Xfanout166 _1060_ VGND VGND VDPWR VDPWR net166 sky130_fd_sc_hd__buf_2
Xfanout100 _1136_ VGND VGND VDPWR VDPWR net100 sky130_fd_sc_hd__buf_4
Xfanout199 net200 VGND VGND VDPWR VDPWR net199 sky130_fd_sc_hd__clkbuf_2
Xfanout122 _1128_ VGND VGND VDPWR VDPWR net122 sky130_fd_sc_hd__buf_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[54\].gen_latches\[4\].p_latch net211 dig_ctrl_inst.latch_mem_inst.gclk\[54\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[54\]\[4\] sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_29_Right_29 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_40_402 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_38_Right_38 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[43\].gen_latches\[2\].p_latch net227 dig_ctrl_inst.latch_mem_inst.gclk\[43\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[43\]\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_20_201 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_234 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[32\].gen_latches\[0\].p_latch net243 dig_ctrl_inst.latch_mem_inst.gclk\[32\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[32\]\[0\] sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_47_Right_47 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_71_593 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1962_ dig_ctrl_inst.latch_mem_inst.RAM\[27\]\[6\] _0130_ _0142_ dig_ctrl_inst.latch_mem_inst.RAM\[42\]\[6\]
+ _0663_ VGND VGND VDPWR VDPWR _0668_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_56_Right_56 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_337 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_315 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_1893_ dig_ctrl_inst.latch_mem_inst.RAM\[2\]\[5\] _1133_ _0129_ dig_ctrl_inst.latch_mem_inst.RAM\[26\]\[5\]
+ VGND VGND VDPWR VDPWR _0600_ sky130_fd_sc_hd__a22o_1
XFILLER_0_11_212 VDPWR VGND VDPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_52 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_2376_ clknet_leaf_4_clk _0003_ net177 VGND VGND VDPWR VDPWR dig_ctrl_inst.spi_receiver_inst.spi_cnt\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_65_Right_65 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_97 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_8
X_2514_ clknet_leaf_9_clk _0111_ net141 VGND VGND VDPWR VDPWR dig_ctrl_inst.cpu_inst.cpu_state\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_2445_ clknet_leaf_11_clk _0053_ net140 VGND VGND VDPWR VDPWR dig_ctrl_inst.cpu_inst.r1\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_75_85 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
X_1258_ net263 dig_ctrl_inst.cpu_inst.r1\[5\] net267 VGND VGND VDPWR VDPWR _1106_
+ sky130_fd_sc_hd__and3b_1
X_1327_ net148 net109 net61 VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.data_we\[18\]
+ sky130_fd_sc_hd__and3_2
X_1189_ net170 VGND VGND VDPWR VDPWR _1037_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_19_281 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_74_Right_74 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_197 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_120 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[20\].gen_latches\[7\].p_latch net185 dig_ctrl_inst.latch_mem_inst.gclk\[20\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[20\]\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_6_250 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_178 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_167 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[58\].gen_latches\[5\].p_latch net205 dig_ctrl_inst.latch_mem_inst.gclk\[58\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[58\]\[5\] sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[47\].gen_latches\[3\].p_latch net220 dig_ctrl_inst.latch_mem_inst.gclk\[47\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[47\]\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_40_307 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_23 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_6
X_2230_ _0747_ _0912_ VGND VGND VDPWR VDPWR _0918_ sky130_fd_sc_hd__nand2_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[36\].gen_latches\[1\].p_latch net236 dig_ctrl_inst.latch_mem_inst.gclk\[36\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[36\]\[1\] sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[2\].gen_latches\[7\].p_latch net186 dig_ctrl_inst.latch_mem_inst.gclk\[2\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[2\]\[7\] sky130_fd_sc_hd__dlxtp_1
X_2161_ _0255_ _0258_ _0254_ VGND VGND VDPWR VDPWR _0852_ sky130_fd_sc_hd__o21a_1
X_2092_ _1014_ _0745_ VGND VGND VDPWR VDPWR _0785_ sky130_fd_sc_hd__or2_2
XFILLER_0_61_98 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_76 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_54 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_101 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_8
X_1945_ dig_ctrl_inst.latch_mem_inst.RAM\[25\]\[6\] net117 net91 net65 VGND VGND VDPWR
+ VDPWR _0651_ sky130_fd_sc_hd__and4_1
XFILLER_0_28_197 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_131 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_16_262 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_315 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_156 VDPWR VGND VDPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_297 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_1876_ dig_ctrl_inst.latch_mem_inst.RAM\[19\]\[5\] net131 net103 net62 VGND VGND
+ VDPWR VDPWR _0583_ sky130_fd_sc_hd__and4_1
X_2359_ dig_ctrl_inst.cpu_inst.port_o\[5\] net372 _0988_ VGND VGND VDPWR VDPWR _0108_
+ sky130_fd_sc_hd__mux2_1
X_2428_ clknet_leaf_9_clk _0036_ net142 VGND VGND VDPWR VDPWR dig_ctrl_inst.cpu_inst.data\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_39_398 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[13\].gen_latches\[6\].p_latch net192 dig_ctrl_inst.latch_mem_inst.gclk\[13\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[13\]\[6\] sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_22_298 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_8_Left_86 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_73_600 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_281 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_46 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_13_243 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1730_ dig_ctrl_inst.latch_mem_inst.RAM\[28\]\[2\] net79 net70 _0120_ dig_ctrl_inst.latch_mem_inst.RAM\[17\]\[2\]
+ VGND VGND VDPWR VDPWR _0440_ sky130_fd_sc_hd__a32o_1
XFILLER_0_40_104 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
X_1592_ dig_ctrl_inst.latch_mem_inst.RAM\[6\]\[0\] net122 _1138_ VGND VGND VDPWR VDPWR
+ _0304_ sky130_fd_sc_hd__and3_2
XFILLER_0_31_79 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
X_1661_ dig_ctrl_inst.latch_mem_inst.RAM\[51\]\[1\] net131 net103 net44 VGND VGND
+ VDPWR VDPWR _0372_ sky130_fd_sc_hd__and4_1
X_2213_ _1125_ _0878_ VGND VGND VDPWR VDPWR _0902_ sky130_fd_sc_hd__or2_1
X_2144_ dig_ctrl_inst.cpu_inst.r0\[1\] _0835_ net41 VGND VGND VDPWR VDPWR _0046_ sky130_fd_sc_hd__mux2_1
XFILLER_0_72_64 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[29\].gen_latches\[0\].p_latch net243 dig_ctrl_inst.latch_mem_inst.gclk\[29\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[29\]\[0\] sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_36_379 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2075_ net163 _0742_ _0744_ VGND VGND VDPWR VDPWR _0768_ sky130_fd_sc_hd__or3_4
X_1928_ dig_ctrl_inst.latch_mem_inst.RAM\[28\]\[6\] net77 net65 VGND VGND VDPWR VDPWR
+ _0634_ sky130_fd_sc_hd__and3_2
X_1859_ net253 _0565_ _0276_ VGND VGND VDPWR VDPWR _0030_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_27_324 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[17\].gen_latches\[7\].p_latch net187 dig_ctrl_inst.latch_mem_inst.gclk\[17\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[17\]\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_62_262 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_224 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_115 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_181 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
Xhold91 dig_ctrl_inst.cpu_inst.r3\[2\] VGND VGND VDPWR VDPWR net373 sky130_fd_sc_hd__dlygate4sd3_1
Xhold80 dig_ctrl_inst.cpu_inst.r2\[1\] VGND VGND VDPWR VDPWR net362 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_9_109 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
X_1713_ _0404_ _0420_ _0421_ _0422_ VGND VGND VDPWR VDPWR _0423_ sky130_fd_sc_hd__or4_1
XFILLER_0_5_337 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_304 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_1575_ _0284_ _0286_ _0285_ VGND VGND VDPWR VDPWR _0287_ sky130_fd_sc_hd__nor3_4
X_1644_ dig_ctrl_inst.latch_mem_inst.RAM\[2\]\[1\] net120 net109 VGND VGND VDPWR VDPWR
+ _0355_ sky130_fd_sc_hd__and3_2
XFILLER_0_67_86 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
Xrebuffer23 net304 VGND VGND VDPWR VDPWR net305 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_49_460 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2127_ _0818_ VGND VGND VDPWR VDPWR _0819_ sky130_fd_sc_hd__inv_2
XFILLER_0_13_3 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_281 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_153 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_2058_ _0743_ _0747_ _0749_ _0746_ VGND VGND VDPWR VDPWR _0751_ sky130_fd_sc_hd__or4b_4
XTAP_TAPCELL_ROW_55_496 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_307 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_1360_ net148 _0137_ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.data_we\[35\]
+ sky130_fd_sc_hd__and2_1
X_1291_ net155 _1135_ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.data_we\[3\]
+ sky130_fd_sc_hd__and2_1
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[10\].clock_gate clknet_leaf_0_clk dig_ctrl_inst.latch_mem_inst.data_we\[10\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.gen_gclk\[10\]._gclk sky130_fd_sc_hd__dlclkp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[62\].gen_latches\[0\].p_latch net244 dig_ctrl_inst.latch_mem_inst.gclk\[62\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[62\]\[0\] sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_46_441 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_218 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
X_1627_ net268 _0338_ _0276_ VGND VGND VDPWR VDPWR _0026_ sky130_fd_sc_hd__mux2_1
X_1489_ net161 dig_ctrl_inst.cpu_inst.data\[1\] _0198_ VGND VGND VDPWR VDPWR _0207_
+ sky130_fd_sc_hd__mux2_1
X_1558_ _0233_ _0172_ VGND VGND VDPWR VDPWR _0271_ sky130_fd_sc_hd__nand2b_1
X_2519__269 VGND VGND VDPWR VDPWR _2519__269/HI net269 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_69_577 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_477 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[50\].gen_latches\[7\].p_latch net183 dig_ctrl_inst.latch_mem_inst.gclk\[50\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[50\]\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_2_3 VDPWR VGND VDPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_335 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_422 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2530_ net276 VGND VGND VDPWR VDPWR uio_out[3] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_21_Left_99 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
Xrebuffer3 net283 VGND VGND VDPWR VDPWR net285 sky130_fd_sc_hd__dlygate4sd1_1
X_2461_ clknet_leaf_3_clk net14 net173 VGND VGND VDPWR VDPWR dig_ctrl_inst.synchronizer_mode_i_inst.pipe\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_2392_ clknet_leaf_4_clk net3 net175 VGND VGND VDPWR VDPWR dig_ctrl_inst.synchronizer_port_i_inst\[0\].pipe\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_1343_ net153 net83 net70 VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.data_we\[26\]
+ sky130_fd_sc_hd__and3_2
X_1412_ _1002_ net180 VGND VGND VDPWR VDPWR _0161_ sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_66_558 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1274_ net267 net264 dig_ctrl_inst.cpu_inst.r3\[4\] VGND VGND VDPWR VDPWR _1122_
+ sky130_fd_sc_hd__and3_2
Xwire36 _0621_ VGND VGND VDPWR VDPWR net36 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_46 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_195 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_16_clk clknet_1_0__leaf_clk VGND VGND VDPWR VDPWR clknet_leaf_16_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_14_243 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
Xfanout178 net180 VGND VGND VDPWR VDPWR net178 sky130_fd_sc_hd__buf_2
Xfanout101 _1136_ VGND VGND VDPWR VDPWR net101 sky130_fd_sc_hd__clkbuf_4
Xfanout145 net146 VGND VGND VDPWR VDPWR net145 sky130_fd_sc_hd__clkbuf_4
Xfanout156 _1097_ VGND VGND VDPWR VDPWR net156 sky130_fd_sc_hd__clkbuf_2
Xfanout189 net190 VGND VGND VDPWR VDPWR net189 sky130_fd_sc_hd__buf_2
Xfanout123 net127 VGND VGND VDPWR VDPWR net123 sky130_fd_sc_hd__buf_2
Xfanout112 net113 VGND VGND VDPWR VDPWR net112 sky130_fd_sc_hd__clkbuf_2
Xfanout167 net168 VGND VGND VDPWR VDPWR net167 sky130_fd_sc_hd__buf_2
XFILLER_0_64_176 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_165 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_403 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[43\].gen_latches\[6\].p_latch net193 dig_ctrl_inst.latch_mem_inst.gclk\[43\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[43\]\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_20_268 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_110 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[32\].gen_latches\[4\].p_latch net211 dig_ctrl_inst.latch_mem_inst.gclk\[32\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[32\]\[4\] sky130_fd_sc_hd__dlxtp_1
X_1961_ dig_ctrl_inst.latch_mem_inst.RAM\[9\]\[6\] _1143_ _0148_ dig_ctrl_inst.latch_mem_inst.RAM\[49\]\[6\]
+ _0660_ VGND VGND VDPWR VDPWR _0667_ sky130_fd_sc_hd__a221o_1
X_1892_ dig_ctrl_inst.latch_mem_inst.RAM\[24\]\[5\] _0127_ _0157_ dig_ctrl_inst.latch_mem_inst.RAM\[60\]\[5\]
+ VGND VGND VDPWR VDPWR _0599_ sky130_fd_sc_hd__a22o_1
X_2513_ clknet_leaf_5_clk _0110_ net179 VGND VGND VDPWR VDPWR net24 sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_5_clk clknet_1_1__leaf_clk VGND VGND VDPWR VDPWR clknet_leaf_5_clk sky130_fd_sc_hd__clkbuf_8
X_2375_ clknet_leaf_5_clk _0002_ net177 VGND VGND VDPWR VDPWR dig_ctrl_inst.spi_receiver_inst.spi_cnt\[0\]
+ sky130_fd_sc_hd__dfrtp_4
X_2444_ clknet_leaf_11_clk _0052_ net142 VGND VGND VDPWR VDPWR dig_ctrl_inst.cpu_inst.r0\[7\]
+ sky130_fd_sc_hd__dfrtp_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[21\].gen_latches\[2\].p_latch net226 dig_ctrl_inst.latch_mem_inst.gclk\[21\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[21\]\[2\] sky130_fd_sc_hd__dlxtp_1
X_1326_ net111 net65 VGND VGND VDPWR VDPWR _0121_ sky130_fd_sc_hd__and2_1
X_1257_ _1010_ _1025_ _1103_ VGND VGND VDPWR VDPWR _1105_ sky130_fd_sc_hd__and3_4
X_1188_ _1018_ _1032_ _1033_ _1034_ _1035_ VGND VGND VDPWR VDPWR _1036_ sky130_fd_sc_hd__o41a_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[59\].gen_latches\[0\].p_latch net244 dig_ctrl_inst.latch_mem_inst.gclk\[59\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[59\]\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_46_165 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[10\].gen_latches\[0\].p_latch net240 dig_ctrl_inst.latch_mem_inst.gclk\[10\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[10\]\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_69_202 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_132 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[47\].gen_latches\[7\].p_latch net189 dig_ctrl_inst.latch_mem_inst.gclk\[47\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[47\]\[7\] sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[3\].gen_latches\[2\].p_latch net231 dig_ctrl_inst.latch_mem_inst.gclk\[3\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[3\]\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_29_57 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
X_2160_ _0845_ _0848_ _0850_ VGND VGND VDPWR VDPWR _0851_ sky130_fd_sc_hd__and3_2
XTAP_TAPCELL_ROW_76_620 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[36\].gen_latches\[5\].p_latch net206 dig_ctrl_inst.latch_mem_inst.gclk\[36\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[36\]\[5\] sky130_fd_sc_hd__dlxtp_1
X_2091_ net161 _0783_ VGND VGND VDPWR VDPWR _0784_ sky130_fd_sc_hd__nand2_1
X_1875_ dig_ctrl_inst.latch_mem_inst.RAM\[7\]\[5\] _1139_ _0579_ _0580_ _0581_ VGND
+ VGND VDPWR VDPWR _0582_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_43_113 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
X_1944_ dig_ctrl_inst.latch_mem_inst.RAM\[63\]\[6\] net104 net81 net45 VGND VGND VDPWR
+ VDPWR _0650_ sky130_fd_sc_hd__and4_1
XFILLER_0_9_12 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_16_263 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[25\].gen_latches\[3\].p_latch net216 dig_ctrl_inst.latch_mem_inst.gclk\[25\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[25\]\[3\] sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_input_latches\[3\].n_latch dig_ctrl_inst.data_out\[3\]
+ clknet_leaf_8_clk VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.wdata\[3\]
+ sky130_fd_sc_hd__dlxtn_1
X_2427_ clknet_leaf_9_clk _0035_ net141 VGND VGND VDPWR VDPWR dig_ctrl_inst.cpu_inst.data\[1\]
+ sky130_fd_sc_hd__dfrtp_2
X_1309_ net155 _1145_ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.data_we\[11\]
+ sky130_fd_sc_hd__and2_1
X_2358_ dig_ctrl_inst.cpu_inst.port_o\[4\] net21 _0988_ VGND VGND VDPWR VDPWR _0107_
+ sky130_fd_sc_hd__mux2_1
X_2289_ _0751_ _0880_ _0877_ VGND VGND VDPWR VDPWR _0971_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_43_3 VDPWR VGND VDPWR VGND sky130_ef_sc_hd__decap_12
Xdig_ctrl_inst.latch_mem_inst.gen_words\[14\].gen_latches\[1\].p_latch net235 dig_ctrl_inst.latch_mem_inst.gclk\[14\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[14\]\[1\] sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_39_399 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_293 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_22_299 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_601 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[7\].gen_latches\[3\].p_latch net222 dig_ctrl_inst.latch_mem_inst.gclk\[7\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[7\]\[3\] sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[15\].clock_gate clknet_leaf_1_clk dig_ctrl_inst.latch_mem_inst.data_we\[15\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.gen_gclk\[15\]._gclk sky130_fd_sc_hd__dlclkp_1
XTAP_TAPCELL_ROW_13_244 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_138 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
X_1660_ dig_ctrl_inst.latch_mem_inst.RAM\[7\]\[1\] net127 net108 net101 VGND VGND
+ VDPWR VDPWR _0371_ sky130_fd_sc_hd__and4_1
X_1591_ dig_ctrl_inst.latch_mem_inst.RAM\[54\]\[0\] net94 net45 VGND VGND VDPWR VDPWR
+ _0303_ sky130_fd_sc_hd__and3_2
XFILLER_0_21_341 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_77 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
X_2212_ _1125_ _0878_ VGND VGND VDPWR VDPWR _0901_ sky130_fd_sc_hd__nand2_1
X_2143_ _0753_ _0830_ _0834_ _0755_ _0833_ VGND VGND VDPWR VDPWR _0835_ sky130_fd_sc_hd__a221o_1
XFILLER_0_72_32 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_208 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[29\].gen_latches\[4\].p_latch net214 dig_ctrl_inst.latch_mem_inst.gclk\[29\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[29\]\[4\] sky130_fd_sc_hd__dlxtp_1
X_2074_ _0264_ _0760_ _0766_ _1068_ VGND VGND VDPWR VDPWR _0767_ sky130_fd_sc_hd__o22a_1
XFILLER_0_8_324 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
XFILLER_0_56_260 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_1858_ _0565_ VGND VGND VDPWR VDPWR _0566_ sky130_fd_sc_hd__inv_2
X_1927_ dig_ctrl_inst.latch_mem_inst.RAM\[39\]\[6\] net103 net99 net55 VGND VGND VDPWR
+ VDPWR _0633_ sky130_fd_sc_hd__and4_1
XFILLER_0_12_330 VDPWR VGND VDPWR VGND sky130_ef_sc_hd__decap_12
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[31\].clock_buffer dig_ctrl_inst.latch_mem_inst.gen_gclk\[31\]._gclk
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.gclk\[31\] sky130_fd_sc_hd__clkbuf_4
X_1789_ dig_ctrl_inst.latch_mem_inst.RAM\[13\]\[3\] _0114_ _0495_ _0496_ _0497_ VGND
+ VGND VDPWR VDPWR _0498_ sky130_fd_sc_hd__a2111o_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[18\].gen_latches\[2\].p_latch net226 dig_ctrl_inst.latch_mem_inst.gclk\[18\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[18\]\[2\] sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_27_325 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_225 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold70 dig_ctrl_inst.cpu_inst.r3\[6\] VGND VGND VDPWR VDPWR net352 sky130_fd_sc_hd__dlygate4sd3_1
Xhold81 dig_ctrl_inst.cpu_inst.r2\[6\] VGND VGND VDPWR VDPWR net363 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_25 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
Xhold92 dig_ctrl_inst.cpu_inst.r1\[0\] VGND VGND VDPWR VDPWR net374 sky130_fd_sc_hd__dlygate4sd3_1
X_1712_ dig_ctrl_inst.latch_mem_inst.RAM\[9\]\[2\] _1143_ _0278_ dig_ctrl_inst.latch_mem_inst.RAM\[5\]\[2\]
+ VGND VGND VDPWR VDPWR _0422_ sky130_fd_sc_hd__a22o_1
XANTENNA_1 _0325_ VGND VGND VDPWR VDPWR sky130_fd_sc_hd__diode_2
X_1643_ dig_ctrl_inst.latch_mem_inst.RAM\[24\]\[1\] net87 net63 VGND VGND VDPWR VDPWR
+ _0354_ sky130_fd_sc_hd__and3_2
X_1574_ _1143_ _1148_ _0116_ _0117_ VGND VGND VDPWR VDPWR _0286_ sky130_fd_sc_hd__or4_4
XFILLER_0_21_193 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_49_461 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer13 _1073_ VGND VGND VDPWR VDPWR net295 sky130_fd_sc_hd__dlygate4sd1_1
X_2126_ _0768_ _0816_ _0817_ _0765_ VGND VGND VDPWR VDPWR _0818_ sky130_fd_sc_hd__o22ai_1
X_2057_ _1011_ net283 VGND VGND VDPWR VDPWR _0750_ sky130_fd_sc_hd__or2_2
XTAP_TAPCELL_ROW_24_306 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_497 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1290_ net132 net126 net106 VGND VGND VDPWR VDPWR _1135_ sky130_fd_sc_hd__and3_4
XTAP_TAPCELL_ROW_46_442 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[62\].gen_latches\[4\].p_latch net214 dig_ctrl_inst.latch_mem_inst.gclk\[62\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[62\]\[4\] sky130_fd_sc_hd__dlxtp_1
X_1626_ _0324_ _0326_ _0337_ _0288_ dig_ctrl_inst.latch_mem_inst.RAM\[0\]\[0\] VGND
+ VGND VDPWR VDPWR _0338_ sky130_fd_sc_hd__o32a_1
XFILLER_0_5_113 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_341 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_69_578 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[51\].gen_latches\[2\].p_latch net229 dig_ctrl_inst.latch_mem_inst.gclk\[51\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[51\]\[2\] sky130_fd_sc_hd__dlxtp_1
X_1488_ _0206_ dig_ctrl_inst.cpu_inst.ip\[0\] _0204_ VGND VGND VDPWR VDPWR _0019_
+ sky130_fd_sc_hd__mux2_1
X_1557_ net138 _0236_ _0167_ VGND VGND VDPWR VDPWR _0270_ sky130_fd_sc_hd__nand3b_1
X_2109_ dig_ctrl_inst.cpu_inst.data\[0\] _0800_ _0801_ VGND VGND VDPWR VDPWR _0802_
+ sky130_fd_sc_hd__and3b_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[40\].gen_latches\[0\].p_latch net244 dig_ctrl_inst.latch_mem_inst.gclk\[40\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[40\]\[0\] sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_52_478 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_185 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_423 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2460_ clknet_leaf_11_clk _0068_ net140 VGND VGND VDPWR VDPWR dig_ctrl_inst.cpu_inst.r2\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_23_288 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
Xrebuffer4 net283 VGND VGND VDPWR VDPWR net286 sky130_fd_sc_hd__dlygate4sd1_1
X_1342_ net83 net69 VGND VGND VDPWR VDPWR _0129_ sky130_fd_sc_hd__and2_2
X_2391_ clknet_leaf_4_clk net342 net179 VGND VGND VDPWR VDPWR dig_ctrl_inst.synchronizer_port_i_inst\[1\].out
+ sky130_fd_sc_hd__dfrtp_1
X_1273_ net263 dig_ctrl_inst.cpu_inst.r1\[4\] net267 VGND VGND VDPWR VDPWR _1121_
+ sky130_fd_sc_hd__and3b_1
X_1411_ net152 _0160_ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.data_we\[63\]
+ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_66_559 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire37 net38 VGND VGND VDPWR VDPWR net37 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_58_174 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[24\].clock_buffer dig_ctrl_inst.latch_mem_inst.gen_gclk\[24\]._gclk
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.gclk\[24\] sky130_fd_sc_hd__clkbuf_4
X_1609_ dig_ctrl_inst.latch_mem_inst.RAM\[46\]\[0\] net72 net58 _0138_ dig_ctrl_inst.latch_mem_inst.RAM\[37\]\[0\]
+ VGND VGND VDPWR VDPWR _0321_ sky130_fd_sc_hd__a32o_1
Xfanout102 net105 VGND VGND VDPWR VDPWR net102 sky130_fd_sc_hd__buf_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[55\].gen_latches\[3\].p_latch net216 dig_ctrl_inst.latch_mem_inst.gclk\[55\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[55\]\[3\] sky130_fd_sc_hd__dlxtp_1
Xfanout179 net180 VGND VGND VDPWR VDPWR net179 sky130_fd_sc_hd__clkbuf_4
Xfanout124 net125 VGND VGND VDPWR VDPWR net124 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_57_504 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout146 net147 VGND VGND VDPWR VDPWR net146 sky130_fd_sc_hd__buf_2
Xfanout135 _1062_ VGND VGND VDPWR VDPWR net135 sky130_fd_sc_hd__buf_4
Xfanout157 net158 VGND VGND VDPWR VDPWR net157 sky130_fd_sc_hd__buf_2
Xfanout168 _1054_ VGND VGND VDPWR VDPWR net168 sky130_fd_sc_hd__dlymetal6s2s_1
X_2532__278 VGND VGND VDPWR VDPWR _2532__278/HI net278 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_40_404 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[44\].gen_latches\[1\].p_latch net234 dig_ctrl_inst.latch_mem_inst.gclk\[44\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[44\]\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_20_247 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_5_192 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1960_ _0656_ _0646_ _0648_ _0644_ VGND VGND VDPWR VDPWR _0666_ sky130_fd_sc_hd__or4_4
XFILLER_0_50_79 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_1891_ _0594_ _0595_ _0596_ _0597_ VGND VGND VDPWR VDPWR _0598_ sky130_fd_sc_hd__or4_1
X_2512_ clknet_leaf_5_clk _0109_ net179 VGND VGND VDPWR VDPWR net23 sky130_fd_sc_hd__dfrtp_1
X_2443_ clknet_leaf_10_clk _0051_ net142 VGND VGND VDPWR VDPWR dig_ctrl_inst.cpu_inst.r0\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_11_225 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[22\].clock_gate clknet_leaf_17_clk dig_ctrl_inst.latch_mem_inst.data_we\[22\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.gen_gclk\[22\]._gclk sky130_fd_sc_hd__dlclkp_1
X_1325_ net155 _0120_ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.data_we\[17\]
+ sky130_fd_sc_hd__and2_1
X_2374_ net282 net2 VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.rst_ni sky130_fd_sc_hd__dfxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[21\].gen_latches\[6\].p_latch net198 dig_ctrl_inst.latch_mem_inst.gclk\[21\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[21\]\[6\] sky130_fd_sc_hd__dlxtp_1
X_1256_ _1103_ VGND VGND VDPWR VDPWR _1104_ sky130_fd_sc_hd__inv_2
X_1187_ net260 net256 dig_ctrl_inst.cpu_inst.r0\[3\] VGND VGND VDPWR VDPWR _1035_
+ sky130_fd_sc_hd__or3_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[59\].gen_latches\[4\].p_latch net214 dig_ctrl_inst.latch_mem_inst.gclk\[59\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[59\]\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_61_169 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_136 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_49_Left_127 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_155 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_339 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_285 VDPWR VGND VDPWR VGND sky130_ef_sc_hd__decap_12
Xdig_ctrl_inst.latch_mem_inst.gen_words\[10\].gen_latches\[4\].p_latch net208 dig_ctrl_inst.latch_mem_inst.gclk\[10\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[10\]\[4\] sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_58_Left_136 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[48\].gen_latches\[2\].p_latch net225 dig_ctrl_inst.latch_mem_inst.gclk\[48\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[48\]\[2\] sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_67_Left_145 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_76_Left_154 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[3\].gen_latches\[6\].p_latch net196 dig_ctrl_inst.latch_mem_inst.gclk\[3\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[3\]\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_60_180 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_136 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[37\].gen_latches\[0\].p_latch net245 dig_ctrl_inst.latch_mem_inst.gclk\[37\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[37\]\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_20_49 VDPWR VGND VDPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_621 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_46 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_8
X_2090_ net254 _1015_ net258 VGND VGND VDPWR VDPWR _0783_ sky130_fd_sc_hd__nor3b_4
XFILLER_0_61_23 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_57 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_15 VDPWR VGND VDPWR VGND sky130_ef_sc_hd__decap_12
X_1943_ dig_ctrl_inst.latch_mem_inst.RAM\[8\]\[6\] net125 net88 VGND VGND VDPWR VDPWR
+ _0649_ sky130_fd_sc_hd__and3_2
X_1874_ dig_ctrl_inst.latch_mem_inst.RAM\[36\]\[5\] net97 net59 VGND VGND VDPWR VDPWR
+ _0581_ sky130_fd_sc_hd__and3_2
XFILLER_0_43_169 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_155 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_8
Xdig_ctrl_inst.latch_mem_inst.gen_input_latches\[7\].n_latch dig_ctrl_inst.data_out\[7\]
+ clknet_leaf_8_clk VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.wdata\[7\]
+ sky130_fd_sc_hd__dlxtn_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[25\].gen_latches\[7\].p_latch net189 dig_ctrl_inst.latch_mem_inst.gclk\[25\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[25\]\[7\] sky130_fd_sc_hd__dlxtp_1
X_2426_ clknet_leaf_8_clk _0034_ net143 VGND VGND VDPWR VDPWR dig_ctrl_inst.cpu_inst.data\[0\]
+ sky130_fd_sc_hd__dfrtp_4
X_2357_ dig_ctrl_inst.cpu_inst.port_o\[3\] net386 _0988_ VGND VGND VDPWR VDPWR _0106_
+ sky130_fd_sc_hd__mux2_1
X_1308_ net106 net126 net92 VGND VGND VDPWR VDPWR _1145_ sky130_fd_sc_hd__and3_4
X_2288_ net369 _0970_ _0967_ VGND VGND VDPWR VDPWR _0055_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_3 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_1239_ net266 net262 dig_ctrl_inst.cpu_inst.r3\[1\] VGND VGND VDPWR VDPWR _1087_
+ sky130_fd_sc_hd__and3_2
XFILLER_0_19_80 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_91 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_125 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[14\].gen_latches\[5\].p_latch net201 dig_ctrl_inst.latch_mem_inst.gclk\[14\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[14\]\[5\] sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_73_602 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[7\].gen_latches\[7\].p_latch net188 dig_ctrl_inst.latch_mem_inst.gclk\[7\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[7\]\[7\] sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_13_245 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_125 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_1590_ dig_ctrl_inst.latch_mem_inst.RAM\[60\]\[0\] net78 net48 VGND VGND VDPWR VDPWR
+ _0302_ sky130_fd_sc_hd__and3_2
XFILLER_0_56_23 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_225 VDPWR VGND VDPWR VGND sky130_ef_sc_hd__decap_12
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[17\].clock_buffer dig_ctrl_inst.latch_mem_inst.gen_gclk\[17\]._gclk
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.gclk\[17\] sky130_fd_sc_hd__clkbuf_4
X_2142_ dig_ctrl_inst.synchronizer_port_i_inst\[1\].out _0802_ _0804_ dig_ctrl_inst.spi_data_o\[1\]
+ VGND VGND VDPWR VDPWR _0834_ sky130_fd_sc_hd__a22o_1
XFILLER_0_56_45 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_2073_ net161 _0759_ VGND VGND VDPWR VDPWR _0766_ sky130_fd_sc_hd__nand2_1
X_2211_ _0788_ _0885_ _0889_ _0899_ VGND VGND VDPWR VDPWR _0900_ sky130_fd_sc_hd__o211a_1
XFILLER_0_8_336 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_6
X_1857_ dig_ctrl_inst.latch_mem_inst.RAM\[0\]\[4\] _0288_ _0519_ _0564_ VGND VGND
+ VDPWR VDPWR _0565_ sky130_fd_sc_hd__o22a_2
X_1788_ dig_ctrl_inst.latch_mem_inst.RAM\[8\]\[3\] net122 net87 VGND VGND VDPWR VDPWR
+ _0497_ sky130_fd_sc_hd__and3_2
X_1926_ dig_ctrl_inst.latch_mem_inst.RAM\[61\]\[6\] net116 net80 net43 VGND VGND VDPWR
+ VDPWR _0632_ sky130_fd_sc_hd__and4_1
XFILLER_0_12_320 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
X_2409_ clknet_leaf_5_clk _0017_ net145 VGND VGND VDPWR VDPWR dig_ctrl_inst.cpu_inst.port_o\[6\]
+ sky130_fd_sc_hd__dfrtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[18\].gen_latches\[6\].p_latch net197 dig_ctrl_inst.latch_mem_inst.gclk\[18\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[18\]\[6\] sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_27_326 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_226 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_180 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_128 VDPWR VGND VDPWR VGND sky130_ef_sc_hd__decap_12
Xhold60 dig_ctrl_inst.synchronizer_port_i_inst\[1\].pipe\[0\] VGND VGND VDPWR VDPWR
+ net342 sky130_fd_sc_hd__dlygate4sd3_1
Xhold71 net24 VGND VGND VDPWR VDPWR net353 sky130_fd_sc_hd__dlygate4sd3_1
Xhold93 dig_ctrl_inst.cpu_inst.r1\[3\] VGND VGND VDPWR VDPWR net375 sky130_fd_sc_hd__dlygate4sd3_1
Xhold82 dig_ctrl_inst.cpu_inst.r3\[7\] VGND VGND VDPWR VDPWR net364 sky130_fd_sc_hd__dlygate4sd3_1
X_1711_ dig_ctrl_inst.latch_mem_inst.RAM\[30\]\[2\] net74 net70 _0142_ dig_ctrl_inst.latch_mem_inst.RAM\[42\]\[2\]
+ VGND VGND VDPWR VDPWR _0421_ sky130_fd_sc_hd__a32o_1
XANTENNA_2 _0443_ VGND VGND VDPWR VDPWR sky130_fd_sc_hd__diode_2
XFILLER_0_53_297 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
X_1642_ dig_ctrl_inst.latch_mem_inst.RAM\[20\]\[1\] net96 net64 VGND VGND VDPWR VDPWR
+ _0353_ sky130_fd_sc_hd__and3_2
XFILLER_0_67_66 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[1\].clock_gate clknet_leaf_19_clk dig_ctrl_inst.latch_mem_inst.data_we\[1\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.gen_gclk\[1\]._gclk sky130_fd_sc_hd__dlclkp_1
X_1573_ net132 net119 _1133_ _1142_ _0277_ VGND VGND VDPWR VDPWR _0285_ sky130_fd_sc_hd__a2111o_1
X_2125_ net157 _0779_ VGND VGND VDPWR VDPWR _0817_ sky130_fd_sc_hd__or2_1
X_2056_ _1011_ net284 VGND VGND VDPWR VDPWR _0749_ sky130_fd_sc_hd__nor2_1
Xrebuffer14 dig_ctrl_inst.cpu_inst.instr\[4\] VGND VGND VDPWR VDPWR net296 sky130_fd_sc_hd__dlygate4sd1_1
XTAP_TAPCELL_ROW_24_307 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1909_ dig_ctrl_inst.latch_mem_inst.RAM\[16\]\[5\] net128 net61 VGND VGND VDPWR VDPWR
+ _0616_ sky130_fd_sc_hd__and3_2
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[27\].clock_gate clknet_leaf_1_clk dig_ctrl_inst.latch_mem_inst.data_we\[27\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.gen_gclk\[27\]._gclk sky130_fd_sc_hd__dlclkp_1
XFILLER_0_53_57 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_46_443 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_337 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_136 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
X_1625_ _0287_ _0320_ _0331_ _0336_ VGND VGND VDPWR VDPWR _0337_ sky130_fd_sc_hd__or4_1
X_1556_ _1119_ net159 _0244_ net160 _1104_ VGND VGND VDPWR VDPWR _0269_ sky130_fd_sc_hd__o32a_1
XTAP_TAPCELL_ROW_69_579 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1487_ _1001_ _0205_ _0173_ VGND VGND VDPWR VDPWR _0206_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_109 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
X_2039_ dig_ctrl_inst.cpu_inst.data\[1\] _0398_ _0741_ VGND VGND VDPWR VDPWR _0035_
+ sky130_fd_sc_hd__mux2_1
X_2108_ dig_ctrl_inst.cpu_inst.data\[3\] dig_ctrl_inst.cpu_inst.data\[2\] VGND VGND
+ VDPWR VDPWR _0801_ sky130_fd_sc_hd__nor2_2
XPHY_EDGE_ROW_30_Left_108 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[51\].gen_latches\[6\].p_latch net192 dig_ctrl_inst.latch_mem_inst.gclk\[51\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[51\]\[6\] sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_52_479 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_275 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[40\].gen_latches\[4\].p_latch net208 dig_ctrl_inst.latch_mem_inst.gclk\[40\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[40\]\[4\] sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_43_424 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1410_ net108 net82 net50 VGND VGND VDPWR VDPWR _0160_ sky130_fd_sc_hd__and3_2
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[63\].clock_buffer dig_ctrl_inst.latch_mem_inst.gen_gclk\[63\]._gclk
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.gclk\[63\] sky130_fd_sc_hd__clkbuf_4
Xrebuffer5 net286 VGND VGND VDPWR VDPWR net287 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_23_223 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_2390_ clknet_leaf_4_clk net4 net175 VGND VGND VDPWR VDPWR dig_ctrl_inst.synchronizer_port_i_inst\[1\].pipe\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_64_45 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_35 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_1272_ _1010_ _1025_ _1118_ VGND VGND VDPWR VDPWR _1120_ sky130_fd_sc_hd__and3_2
X_1341_ net148 _0128_ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.data_we\[25\]
+ sky130_fd_sc_hd__and2_1
Xwire38 _0578_ VGND VGND VDPWR VDPWR net38 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_82 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
Xfanout125 net127 VGND VGND VDPWR VDPWR net125 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_66_3 VDPWR VGND VDPWR VGND sky130_ef_sc_hd__decap_12
Xfanout147 dig_ctrl_inst.cpu_inst.rst_ni VGND VGND VDPWR VDPWR net147 sky130_fd_sc_hd__clkbuf_2
X_1608_ dig_ctrl_inst.latch_mem_inst.RAM\[8\]\[0\] _1142_ _0153_ dig_ctrl_inst.latch_mem_inst.RAM\[55\]\[0\]
+ _0319_ VGND VGND VDPWR VDPWR _0320_ sky130_fd_sc_hd__a221o_1
X_1539_ _0249_ _0251_ VGND VGND VDPWR VDPWR _0252_ sky130_fd_sc_hd__nand2_1
Xfanout114 net115 VGND VGND VDPWR VDPWR net114 sky130_fd_sc_hd__buf_4
Xfanout103 net105 VGND VGND VDPWR VDPWR net103 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_57_505 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout169 _1045_ VGND VGND VDPWR VDPWR net169 sky130_fd_sc_hd__buf_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[55\].gen_latches\[7\].p_latch net184 dig_ctrl_inst.latch_mem_inst.gclk\[55\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[55\]\[7\] sky130_fd_sc_hd__dlxtp_1
Xfanout158 _1067_ VGND VGND VDPWR VDPWR net158 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_64_112 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_175 VDPWR VGND VDPWR VGND sky130_ef_sc_hd__decap_12
Xdig_ctrl_inst.latch_mem_inst.gen_words\[0\].gen_latches\[0\].p_latch net246 dig_ctrl_inst.latch_mem_inst.gclk\[0\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[0\]\[0\] sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_40_405 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_337 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[44\].gen_latches\[5\].p_latch net200 dig_ctrl_inst.latch_mem_inst.gclk\[44\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[44\]\[5\] sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[33\].gen_latches\[3\].p_latch net215 dig_ctrl_inst.latch_mem_inst.gclk\[33\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[33\]\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_18_27 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_5_193 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_16_Right_16 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XFILLER_0_70_126 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_134 VDPWR VGND VDPWR VGND sky130_ef_sc_hd__decap_12
X_1890_ dig_ctrl_inst.latch_mem_inst.RAM\[28\]\[5\] net77 net64 _0154_ dig_ctrl_inst.latch_mem_inst.RAM\[57\]\[5\]
+ VGND VGND VDPWR VDPWR _0597_ sky130_fd_sc_hd__a32o_1
XPHY_EDGE_ROW_25_Right_25 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[22\].gen_latches\[1\].p_latch net236 dig_ctrl_inst.latch_mem_inst.gclk\[22\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[22\]\[1\] sky130_fd_sc_hd__dlxtp_1
X_2511_ clknet_leaf_5_clk _0108_ net179 VGND VGND VDPWR VDPWR net22 sky130_fd_sc_hd__dfrtp_1
X_2442_ clknet_leaf_6_clk _0050_ net145 VGND VGND VDPWR VDPWR dig_ctrl_inst.cpu_inst.r0\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_2373_ _0990_ _0996_ _0201_ VGND VGND VDPWR VDPWR _0113_ sky130_fd_sc_hd__o21a_1
X_1324_ net132 net119 net71 VGND VGND VDPWR VDPWR _0120_ sky130_fd_sc_hd__and3_4
X_1186_ net260 dig_ctrl_inst.cpu_inst.r2\[3\] VGND VGND VDPWR VDPWR _1034_ sky130_fd_sc_hd__and2b_1
X_1255_ _1018_ _1099_ _1100_ _1101_ _1102_ VGND VGND VDPWR VDPWR _1103_ sky130_fd_sc_hd__o41a_4
XPHY_EDGE_ROW_34_Right_34 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_315 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_337 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_43_Right_43 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_340 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_253 VDPWR VGND VDPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_297 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_52_Right_52 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[4\].gen_latches\[1\].p_latch net237 dig_ctrl_inst.latch_mem_inst.gclk\[4\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[4\]\[1\] sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_2_174 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[48\].gen_latches\[6\].p_latch net192 dig_ctrl_inst.latch_mem_inst.gclk\[48\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[48\]\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_77_281 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_61_Right_61 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_148 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_189 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_70_Right_70 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[37\].gen_latches\[4\].p_latch net208 dig_ctrl_inst.latch_mem_inst.gclk\[37\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[37\]\[4\] sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_76_622 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[6\].clock_gate clknet_leaf_17_clk dig_ctrl_inst.latch_mem_inst.data_we\[6\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.gen_gclk\[6\]._gclk sky130_fd_sc_hd__dlclkp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[26\].gen_latches\[2\].p_latch net230 dig_ctrl_inst.latch_mem_inst.gclk\[26\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[26\]\[2\] sky130_fd_sc_hd__dlxtp_1
X_1942_ dig_ctrl_inst.latch_mem_inst.RAM\[3\]\[6\] net132 net124 net107 VGND VGND
+ VDPWR VDPWR _0648_ sky130_fd_sc_hd__and4_1
XFILLER_0_61_57 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_123 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_27 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_1873_ dig_ctrl_inst.latch_mem_inst.RAM\[39\]\[5\] net107 net101 net59 VGND VGND
+ VDPWR VDPWR _0580_ sky130_fd_sc_hd__and4_1
XFILLER_0_43_126 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_178 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_278 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
X_2356_ dig_ctrl_inst.cpu_inst.port_o\[2\] net385 _0988_ VGND VGND VDPWR VDPWR _0105_
+ sky130_fd_sc_hd__mux2_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[15\].gen_latches\[0\].p_latch net243 dig_ctrl_inst.latch_mem_inst.gclk\[15\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[15\]\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_10_83 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_2425_ clknet_leaf_13_clk _0033_ net139 VGND VGND VDPWR VDPWR dig_ctrl_inst.cpu_inst.instr\[7\]
+ sky130_fd_sc_hd__dfrtp_2
X_1307_ net154 net124 net83 VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.data_we\[10\]
+ sky130_fd_sc_hd__and3_2
X_2287_ _0751_ _0856_ _0854_ VGND VGND VDPWR VDPWR _0970_ sky130_fd_sc_hd__o21ai_1
X_1238_ net262 dig_ctrl_inst.cpu_inst.r1\[1\] net266 VGND VGND VDPWR VDPWR _1086_
+ sky130_fd_sc_hd__and3b_1
XFILLER_0_29_3 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_8
X_1169_ dig_ctrl_inst.cpu_inst.instr\[7\] net253 dig_ctrl_inst.cpu_inst.instr\[6\]
+ net252 VGND VGND VDPWR VDPWR _1017_ sky130_fd_sc_hd__or4_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[8\].gen_latches\[2\].p_latch net225 dig_ctrl_inst.latch_mem_inst.gclk\[8\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[8\]\[2\] sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_73_603 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_390 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_17 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[56\].clock_buffer dig_ctrl_inst.latch_mem_inst.gen_gclk\[56\]._gclk
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.gclk\[56\] sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_21_290 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_204 VDPWR VGND VDPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_237 VDPWR VGND VDPWR VGND sky130_ef_sc_hd__decap_12
X_2210_ _0750_ _0892_ _0893_ _0898_ VGND VGND VDPWR VDPWR _0899_ sky130_fd_sc_hd__o211a_1
XFILLER_0_72_12 VDPWR VGND VDPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_57 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
X_2141_ _0820_ _0822_ _0832_ VGND VGND VDPWR VDPWR _0833_ sky130_fd_sc_hd__nand3_1
X_2072_ net163 _0764_ VGND VGND VDPWR VDPWR _0765_ sky130_fd_sc_hd__nand2_2
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[34\].clock_gate clknet_leaf_17_clk dig_ctrl_inst.latch_mem_inst.data_we\[34\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.gen_gclk\[34\]._gclk sky130_fd_sc_hd__dlclkp_1
XFILLER_0_8_315 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_1925_ dig_ctrl_inst.latch_mem_inst.RAM\[50\]\[6\] net110 net43 VGND VGND VDPWR VDPWR
+ _0631_ sky130_fd_sc_hd__and3_2
X_1856_ _0534_ _0551_ _0558_ _0563_ VGND VGND VDPWR VDPWR _0564_ sky130_fd_sc_hd__or4_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[19\].gen_latches\[1\].p_latch net239 dig_ctrl_inst.latch_mem_inst.gclk\[19\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[19\]\[1\] sky130_fd_sc_hd__dlxtp_1
X_1787_ dig_ctrl_inst.latch_mem_inst.RAM\[43\]\[3\] net104 net91 net56 VGND VGND VDPWR
+ VDPWR _0496_ sky130_fd_sc_hd__and4_1
X_2339_ dig_ctrl_inst.cpu_inst.port_o\[3\] dig_ctrl_inst.spi_data_i\[3\] _0986_ VGND
+ VGND VDPWR VDPWR _0090_ sky130_fd_sc_hd__mux2_1
X_2408_ clknet_leaf_6_clk _0016_ net145 VGND VGND VDPWR VDPWR dig_ctrl_inst.cpu_inst.port_o\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_2_Right_2 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_27_327 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_232 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_10_227 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold50 dig_ctrl_inst.synchronizer_port_i_inst\[4\].pipe\[0\] VGND VGND VDPWR VDPWR
+ net332 sky130_fd_sc_hd__dlygate4sd3_1
Xhold94 dig_ctrl_inst.cpu_inst.r3\[4\] VGND VGND VDPWR VDPWR net376 sky130_fd_sc_hd__dlygate4sd3_1
Xhold61 dig_ctrl_inst.stb_d VGND VGND VDPWR VDPWR net343 sky130_fd_sc_hd__dlygate4sd3_1
Xhold83 dig_ctrl_inst.cpu_inst.r1\[5\] VGND VGND VDPWR VDPWR net365 sky130_fd_sc_hd__dlygate4sd3_1
Xhold72 dig_ctrl_inst.cpu_inst.prev_state\[2\] VGND VGND VDPWR VDPWR net354 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_295 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_251 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_1572_ _0280_ _0281_ _0282_ _0283_ VGND VGND VDPWR VDPWR _0284_ sky130_fd_sc_hd__or4_2
X_1710_ dig_ctrl_inst.latch_mem_inst.RAM\[21\]\[2\] _0124_ _0151_ dig_ctrl_inst.latch_mem_inst.RAM\[53\]\[2\]
+ _0415_ VGND VGND VDPWR VDPWR _0420_ sky130_fd_sc_hd__a221o_1
XANTENNA_3 _0477_ VGND VGND VDPWR VDPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_26 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
X_1641_ dig_ctrl_inst.latch_mem_inst.RAM\[21\]\[1\] net116 net99 net62 VGND VGND VDPWR
+ VDPWR _0352_ sky130_fd_sc_hd__and4_1
XFILLER_0_6_48 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
X_2124_ _0814_ _0815_ VGND VGND VDPWR VDPWR _0816_ sky130_fd_sc_hd__nor2_1
Xrebuffer15 _1026_ VGND VGND VDPWR VDPWR net297 sky130_fd_sc_hd__buf_6
XFILLER_0_8_101 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
X_2055_ _1015_ _1031_ VGND VGND VDPWR VDPWR _0748_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_24_308 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1839_ dig_ctrl_inst.latch_mem_inst.RAM\[34\]\[4\] net111 net58 VGND VGND VDPWR VDPWR
+ _0547_ sky130_fd_sc_hd__and3_2
XFILLER_0_32_70 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_295 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_340 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
X_1908_ dig_ctrl_inst.latch_mem_inst.RAM\[61\]\[5\] _0158_ _0612_ _0613_ _0614_ VGND
+ VGND VDPWR VDPWR _0615_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_12_29 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[63\].gen_latches\[3\].p_latch net220 dig_ctrl_inst.latch_mem_inst.gclk\[63\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[63\]\[3\] sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[52\].gen_latches\[1\].p_latch net239 dig_ctrl_inst.latch_mem_inst.gclk\[52\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[52\]\[1\] sky130_fd_sc_hd__dlxtp_1
X_1624_ _0332_ _0333_ _0334_ _0335_ VGND VGND VDPWR VDPWR _0336_ sky130_fd_sc_hd__or4_1
X_1555_ _0245_ _0267_ VGND VGND VDPWR VDPWR _0268_ sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_19_clk clknet_1_1__leaf_clk VGND VGND VDPWR VDPWR clknet_leaf_19_clk
+ sky130_fd_sc_hd__clkbuf_8
X_2107_ dig_ctrl_inst.cpu_inst.data\[1\] _0799_ VGND VGND VDPWR VDPWR _0800_ sky130_fd_sc_hd__nor2_1
X_1486_ net164 dig_ctrl_inst.cpu_inst.data\[0\] _0198_ VGND VGND VDPWR VDPWR _0205_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_313 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
X_2038_ dig_ctrl_inst.cpu_inst.data\[0\] _0338_ _0741_ VGND VGND VDPWR VDPWR _0034_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_3 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_221 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_192 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[49\].clock_buffer dig_ctrl_inst.latch_mem_inst.gen_gclk\[49\]._gclk
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.gclk\[49\] sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_43_425 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_25 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
Xrebuffer6 net287 VGND VGND VDPWR VDPWR net288 sky130_fd_sc_hd__dlygate4sd1_1
X_1340_ net114 net90 net61 VGND VGND VDPWR VDPWR _0128_ sky130_fd_sc_hd__and3_2
X_1271_ _1118_ VGND VGND VDPWR VDPWR _1119_ sky130_fd_sc_hd__inv_2
Xwire39 net40 VGND VGND VDPWR VDPWR net39 sky130_fd_sc_hd__clkbuf_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[56\].gen_latches\[2\].p_latch net229 dig_ctrl_inst.latch_mem_inst.gclk\[56\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[56\]\[2\] sky130_fd_sc_hd__dlxtp_1
Xclkbuf_leaf_8_clk clknet_1_1__leaf_clk VGND VGND VDPWR VDPWR clknet_leaf_8_clk sky130_fd_sc_hd__clkbuf_8
X_1469_ _0195_ dig_ctrl_inst.spi_addr\[5\] _0186_ VGND VGND VDPWR VDPWR _0197_ sky130_fd_sc_hd__or3b_1
Xfanout126 net127 VGND VGND VDPWR VDPWR net126 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_59_3 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_80 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
Xfanout104 net105 VGND VGND VDPWR VDPWR net104 sky130_fd_sc_hd__buf_2
X_1538_ net170 net169 VGND VGND VDPWR VDPWR _0251_ sky130_fd_sc_hd__or2_1
Xfanout148 net151 VGND VGND VDPWR VDPWR net148 sky130_fd_sc_hd__clkbuf_2
Xfanout115 net116 VGND VGND VDPWR VDPWR net115 sky130_fd_sc_hd__buf_4
X_1607_ dig_ctrl_inst.latch_mem_inst.RAM\[51\]\[0\] _0149_ _0150_ dig_ctrl_inst.latch_mem_inst.RAM\[52\]\[0\]
+ VGND VGND VDPWR VDPWR _0319_ sky130_fd_sc_hd__a22o_1
Xfanout159 _1125_ VGND VGND VDPWR VDPWR net159 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_57_506 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[45\].gen_latches\[0\].p_latch net243 dig_ctrl_inst.latch_mem_inst.gclk\[45\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[45\]\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_49_187 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_40_406 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[0\].gen_latches\[4\].p_latch net211 dig_ctrl_inst.latch_mem_inst.gclk\[0\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[0\]\[4\] sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_5_194 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_3 VDPWR VGND VDPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_113 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[33\].gen_latches\[7\].p_latch net183 dig_ctrl_inst.latch_mem_inst.gclk\[33\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[33\]\[7\] sky130_fd_sc_hd__dlxtp_1
X_2510_ clknet_leaf_5_clk _0107_ net179 VGND VGND VDPWR VDPWR net21 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_149 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[39\].clock_gate clknet_leaf_2_clk dig_ctrl_inst.latch_mem_inst.data_we\[39\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.gen_gclk\[39\]._gclk sky130_fd_sc_hd__dlclkp_1
XFILLER_0_55_146 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_341 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_59 VDPWR VGND VDPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_48 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
XFILLER_0_59_79 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_2441_ clknet_leaf_6_clk _0049_ net145 VGND VGND VDPWR VDPWR dig_ctrl_inst.cpu_inst.r0\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_2372_ _1027_ dig_ctrl_inst.cpu_inst.cpu_state\[1\] _0990_ VGND VGND VDPWR VDPWR
+ _0112_ sky130_fd_sc_hd__mux2_1
X_1323_ net128 net150 net62 VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.data_we\[16\]
+ sky130_fd_sc_hd__and3_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[22\].gen_latches\[5\].p_latch net200 dig_ctrl_inst.latch_mem_inst.gclk\[22\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[22\]\[5\] sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[11\].gen_latches\[3\].p_latch net222 dig_ctrl_inst.latch_mem_inst.gclk\[11\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[11\]\[3\] sky130_fd_sc_hd__dlxtp_1
X_1185_ net257 dig_ctrl_inst.cpu_inst.r1\[3\] VGND VGND VDPWR VDPWR _1033_ sky130_fd_sc_hd__and2b_1
X_1254_ net260 net257 dig_ctrl_inst.cpu_inst.r0\[5\] VGND VGND VDPWR VDPWR _1102_
+ sky130_fd_sc_hd__or3_1
XFILLER_0_6_243 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[49\].gen_latches\[1\].p_latch net237 dig_ctrl_inst.latch_mem_inst.gclk\[49\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[49\]\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_6_265 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_8
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[20\].clock_buffer dig_ctrl_inst.latch_mem_inst.gen_gclk\[20\]._gclk
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.gclk\[20\] sky130_fd_sc_hd__clkbuf_4
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[6\].clock_buffer dig_ctrl_inst.latch_mem_inst.gen_gclk\[6\]._gclk
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.gclk\[6\] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_4_81 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_260 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[41\].clock_gate clknet_leaf_13_clk dig_ctrl_inst.latch_mem_inst.data_we\[41\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.gen_gclk\[41\]._gclk sky130_fd_sc_hd__dlclkp_1
XFILLER_0_37_113 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_175 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[4\].gen_latches\[5\].p_latch net204 dig_ctrl_inst.latch_mem_inst.gclk\[4\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[4\]\[5\] sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_76_623 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1872_ dig_ctrl_inst.latch_mem_inst.RAM\[42\]\[5\] net83 net59 VGND VGND VDPWR VDPWR
+ _0579_ sky130_fd_sc_hd__and3_2
X_1941_ dig_ctrl_inst.latch_mem_inst.RAM\[59\]\[6\] net107 net92 net48 VGND VGND VDPWR
+ VDPWR _0647_ sky130_fd_sc_hd__and4_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[26\].gen_latches\[6\].p_latch net194 dig_ctrl_inst.latch_mem_inst.gclk\[26\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[26\]\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_3_213 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[15\].gen_latches\[4\].p_latch net214 dig_ctrl_inst.latch_mem_inst.gclk\[15\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[15\]\[4\] sky130_fd_sc_hd__dlxtp_1
X_2355_ dig_ctrl_inst.cpu_inst.port_o\[1\] net392 _0988_ VGND VGND VDPWR VDPWR _0104_
+ sky130_fd_sc_hd__mux2_1
X_1306_ net290 _1078_ net134 _1062_ net136 VGND VGND VDPWR VDPWR _1144_ sky130_fd_sc_hd__a2111oi_4
X_2286_ net367 _0969_ _0967_ VGND VGND VDPWR VDPWR _0054_ sky130_fd_sc_hd__mux2_1
X_2424_ clknet_leaf_13_clk _0032_ net139 VGND VGND VDPWR VDPWR dig_ctrl_inst.cpu_inst.instr\[6\]
+ sky130_fd_sc_hd__dfrtp_2
X_1237_ _1010_ _1025_ net163 VGND VGND VDPWR VDPWR _1085_ sky130_fd_sc_hd__and3_2
X_1168_ net252 net253 VGND VGND VDPWR VDPWR _1016_ sky130_fd_sc_hd__or2_1
XFILLER_0_19_113 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
XFILLER_0_59_293 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_341 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_73_604 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[8\].gen_latches\[6\].p_latch net196 dig_ctrl_inst.latch_mem_inst.gclk\[8\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[8\]\[6\] sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_38_391 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_17 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_216 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_21_291 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_138 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_249 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
X_2140_ _0257_ _0787_ _0824_ _0827_ _0831_ VGND VGND VDPWR VDPWR _0832_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_72_24 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
X_2071_ _0742_ _0744_ VGND VGND VDPWR VDPWR _0764_ sky130_fd_sc_hd__nor2_1
X_1924_ dig_ctrl_inst.latch_mem_inst.RAM\[58\]\[6\] net84 net50 VGND VGND VDPWR VDPWR
+ _0630_ sky130_fd_sc_hd__and3_2
X_1855_ _0559_ _0560_ _0561_ _0562_ VGND VGND VDPWR VDPWR _0563_ sky130_fd_sc_hd__or4_1
XFILLER_0_16_116 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_138 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
X_1786_ dig_ctrl_inst.latch_mem_inst.RAM\[29\]\[3\] net119 net82 net71 VGND VGND VDPWR
+ VDPWR _0495_ sky130_fd_sc_hd__and4_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[19\].gen_latches\[5\].p_latch net200 dig_ctrl_inst.latch_mem_inst.gclk\[19\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[19\]\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_12_300 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_8
X_2338_ dig_ctrl_inst.cpu_inst.port_o\[2\] dig_ctrl_inst.spi_data_i\[2\] _0986_ VGND
+ VGND VDPWR VDPWR _0089_ sky130_fd_sc_hd__mux2_1
X_2407_ clknet_leaf_6_clk _0015_ net145 VGND VGND VDPWR VDPWR dig_ctrl_inst.cpu_inst.port_o\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_41_3 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_6
X_2269_ net167 _0860_ _0954_ net170 VGND VGND VDPWR VDPWR _0955_ sky130_fd_sc_hd__a211o_1
XFILLER_0_39_208 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_35_372 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_328 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_82 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_4
Xhold40 dig_ctrl_inst.latch_mem_inst.wdata\[6\] VGND VGND VDPWR VDPWR net322 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_174 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
Xhold62 dig_ctrl_inst.spi_receiver_inst.spi_sclk_sync VGND VGND VDPWR VDPWR net344
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold73 dig_ctrl_inst.spi_miso_o VGND VGND VDPWR VDPWR net355 sky130_fd_sc_hd__dlygate4sd3_1
Xhold51 dig_ctrl_inst.spi_receiver_inst.synchronizer_spi_sclk.pipe\[0\] VGND VGND
+ VDPWR VDPWR net333 sky130_fd_sc_hd__dlygate4sd3_1
Xhold84 dig_ctrl_inst.cpu_inst.r2\[5\] VGND VGND VDPWR VDPWR net366 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_16 VDPWR VGND VDPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_39 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
Xhold95 dig_ctrl_inst.cpu_inst.r1\[7\] VGND VGND VDPWR VDPWR net377 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_49 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_6
X_1571_ _1093_ net123 net92 VGND VGND VDPWR VDPWR _0283_ sky130_fd_sc_hd__and3_2
XANTENNA_4 _0511_ VGND VGND VDPWR VDPWR sky130_fd_sc_hd__diode_2
XFILLER_0_21_185 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
X_1640_ dig_ctrl_inst.latch_mem_inst.RAM\[47\]\[1\] net104 net81 net56 VGND VGND VDPWR
+ VDPWR _0351_ sky130_fd_sc_hd__and4_1
XFILLER_0_67_79 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
Xrebuffer16 net181 VGND VGND VDPWR VDPWR net298 sky130_fd_sc_hd__dlymetal6s2s_1
X_2123_ net157 _0775_ VGND VGND VDPWR VDPWR _0815_ sky130_fd_sc_hd__nor2_1
XFILLER_0_16_83 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
X_2054_ _1015_ _1031_ VGND VGND VDPWR VDPWR _0747_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_24_309 VGND VDPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[13\].clock_buffer dig_ctrl_inst.latch_mem_inst.gen_gclk\[13\]._gclk
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.gclk\[13\] sky130_fd_sc_hd__clkbuf_4
X_1838_ dig_ctrl_inst.latch_mem_inst.RAM\[39\]\[4\] _0139_ _0543_ _0544_ _0545_ VGND
+ VGND VDPWR VDPWR _0546_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_32_82 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_2
X_1907_ dig_ctrl_inst.latch_mem_inst.RAM\[12\]\[5\] net120 net76 VGND VGND VDPWR VDPWR
+ _0614_ sky130_fd_sc_hd__and3_2
X_1769_ dig_ctrl_inst.latch_mem_inst.RAM\[48\]\[3\] net128 net44 VGND VGND VDPWR VDPWR
+ _0478_ sky130_fd_sc_hd__and3_2
XFILLER_0_12_141 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__fill_1
Xoutput30 net30 VGND VGND VDPWR VDPWR uo_out[2] sky130_fd_sc_hd__buf_2
XFILLER_0_35_277 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_16 VGND VGND VDPWR VDPWR sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[63\].gen_latches\[7\].p_latch net185 dig_ctrl_inst.latch_mem_inst.gclk\[63\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[63\]\[7\] sky130_fd_sc_hd__dlxtp_1
X_1623_ dig_ctrl_inst.latch_mem_inst.RAM\[7\]\[0\] _1139_ _0290_ _0300_ _0301_ VGND
+ VGND VDPWR VDPWR _0335_ sky130_fd_sc_hd__a2111o_1
X_1485_ _1030_ _0199_ _0203_ _0201_ VGND VGND VDPWR VDPWR _0204_ sky130_fd_sc_hd__or4b_4
X_1554_ _1037_ net169 _0253_ _0265_ _0266_ VGND VGND VDPWR VDPWR _0267_ sky130_fd_sc_hd__o221a_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[52\].gen_latches\[5\].p_latch net201 dig_ctrl_inst.latch_mem_inst.gclk\[52\]
+ VGND VGND VDPWR VDPWR dig_ctrl_inst.latch_mem_inst.RAM\[52\]\[5\] sky130_fd_sc_hd__dlxtp_1
.ends

